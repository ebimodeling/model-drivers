netcdf all_bced_1960_1999_hadgem2-es_rcp6p0_2005-2099 {
dimensions:
	lat = UNLIMITED ; // (360 currently)
	lon = 720 ;
	time = 34698 ;
variables:
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
	float psAdjust(lat, lon, time) ;
		psAdjust:_FillValue = 1.e+20f ;
		psAdjust:long_name = "Bias-Corrected Sea Level Pressure" ;
		psAdjust:units = "Pa" ;
		psAdjust:standard_name = "air_pressure_at_sea_level" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:units = "days since 1860-01-01 00:00:00" ;
		time:calendar = "standard" ;
	float rldsAdjust(lat, lon, time) ;
		rldsAdjust:_FillValue = 1.e+20f ;
		rldsAdjust:long_name = "Bias-Corrected Surface Downwelling Longwave Radiation" ;
		rldsAdjust:units = "W m-2" ;
		rldsAdjust:standard_name = "surface_downwelling_longwave_flux_in_air" ;
	float rsdsAdjust(lat, lon, time) ;
		rsdsAdjust:_FillValue = 1.e+20f ;
		rsdsAdjust:long_name = "Bias-Corrected Surface Downwelling Shortwave Radiation" ;
		rsdsAdjust:units = "W m-2" ;
		rsdsAdjust:standard_name = "surface_downwelling_shortwave_flux_in_air" ;
	float tasAdjust(lat, lon, time) ;
		tasAdjust:_FillValue = 1.e+20f ;
	float tasmaxAdjust(lat, lon, time) ;
		tasmaxAdjust:_FillValue = 1.e+20f ;
	float tasminAdjust(lat, lon, time) ;
		tasminAdjust:_FillValue = 1.e+20f ;
	float uasAdjust(lat, lon, time) ;
		uasAdjust:_FillValue = 1.e+20f ;
		uasAdjust:long_name = "Bias-Corrected Eastward Near-Surface Wind" ;
		uasAdjust:units = "m s-1" ;
		uasAdjust:standard_name = "eastward_wind" ;
	float vasAdjust(lat, lon, time) ;
		vasAdjust:_FillValue = 1.e+20f ;
		vasAdjust:long_name = "Bias-Corrected Northward Near-Surface Wind" ;
		vasAdjust:units = "m s-1" ;
		vasAdjust:standard_name = "northward_wind" ;
	float prAdjust(lat, lon, time) ;
		prAdjust:_FillValue = 1.e+20f ;
		prAdjust:comment = "includes all types (rain, snow, large-scale, convective, etc.)" ;
		prAdjust:long_name = "Bias-Corrected Precipitation" ;
		prAdjust:units = "kg m-2 s-1" ;
		prAdjust:standard_name = "precipitation_flux" ;

// global attributes:
		:history = "Thu May  8 12:32:15 2014: ncks --no_tmp_fl -A -v Adjust$ pr_bced_1960_1999_hadgem2-es_rcp6p0_2005-2099p.nc all_1960_1999_hadgem2-es_rcp6p0_2005-2099.nc\nThu May  8 12:14:02 2014: ncks --no_tmp_fl -A -v Adjust$ vas_bced_1960_1999_hadgem2-es_rcp6p0_2005-2099p.nc all_1960_1999_hadgem2-es_rcp6p0_2005-2099.nc\nThu May  8 12:00:41 2014: ncks --no_tmp_fl -A -v Adjust$ uas_bced_1960_1999_hadgem2-es_rcp6p0_2005-2099p.nc all_1960_1999_hadgem2-es_rcp6p0_2005-2099.nc\nThu May  8 11:45:54 2014: ncks --no_tmp_fl -A -v Adjust$ tasmin_bced_1960_1999_hadgem2-es_rcp6p0_2005-2099pt.nc all_1960_1999_hadgem2-es_rcp6p0_2005-2099.nc\nThu May  8 11:31:09 2014: ncks --no_tmp_fl -A -v Adjust$ tasmax_bced_1960_1999_hadgem2-es_rcp6p0_2005-2099pt.nc all_1960_1999_hadgem2-es_rcp6p0_2005-2099.nc\nThu May  8 11:16:46 2014: ncks --no_tmp_fl -A -v Adjust$ tas_bced_1960_1999_hadgem2-es_rcp6p0_2005-2099pt.nc all_1960_1999_hadgem2-es_rcp6p0_2005-2099.nc\nThu May  8 11:04:36 2014: ncks --no_tmp_fl -A -v Adjust$ rsds_bced_1960_1999_hadgem2-es_rcp6p0_2005-2099p.nc all_1960_1999_hadgem2-es_rcp6p0_2005-2099.nc\nThu May  8 10:52:14 2014: ncks --no_tmp_fl -A -v Adjust$ rlds_bced_1960_1999_hadgem2-es_rcp6p0_2005-2099p.nc all_1960_1999_hadgem2-es_rcp6p0_2005-2099.nc\nThu May  8 10:40:40 2014: ncks --no_tmp_fl -A -v Adjust$ ps_bced_1960_1999_hadgem2-es_rcp6p0_2005-2099p.nc all_1960_1999_hadgem2-es_rcp6p0_2005-2099.nc" ;
		:NCO = "4.4.2" ;
data:

 time = 52961, 52962, 52963, 52964, 52965, 52966, 52967, 52968, 52969, 52970, 
    52971, 52972, 52973, 52974, 52975, 52976, 52977, 52978, 52979, 52980, 
    52981, 52982, 52983, 52984, 52985, 52986, 52987, 52988, 52989, 52990, 
    52991, 52992, 52993, 52994, 52995, 52996, 52997, 52998, 52999, 53000, 
    53001, 53002, 53003, 53004, 53005, 53006, 53007, 53008, 53009, 53010, 
    53011, 53012, 53013, 53014, 53015, 53016, 53017, 53018, 53019, 53020, 
    53021, 53022, 53023, 53024, 53025, 53026, 53027, 53028, 53029, 53030, 
    53031, 53032, 53033, 53034, 53035, 53036, 53037, 53038, 53039, 53040, 
    53041, 53042, 53043, 53044, 53045, 53046, 53047, 53048, 53049, 53050, 
    53051, 53052, 53053, 53054, 53055, 53056, 53057, 53058, 53059, 53060, 
    53061, 53062, 53063, 53064, 53065, 53066, 53067, 53068, 53069, 53070, 
    53071, 53072, 53073, 53074, 53075, 53076, 53077, 53078, 53079, 53080, 
    53081, 53082, 53083, 53084, 53085, 53086, 53087, 53088, 53089, 53090, 
    53091, 53092, 53093, 53094, 53095, 53096, 53097, 53098, 53099, 53100, 
    53101, 53102, 53103, 53104, 53105, 53106, 53107, 53108, 53109, 53110, 
    53111, 53112, 53113, 53114, 53115, 53116, 53117, 53118, 53119, 53120, 
    53121, 53122, 53123, 53124, 53125, 53126, 53127, 53128, 53129, 53130, 
    53131, 53132, 53133, 53134, 53135, 53136, 53137, 53138, 53139, 53140, 
    53141, 53142, 53143, 53144, 53145, 53146, 53147, 53148, 53149, 53150, 
    53151, 53152, 53153, 53154, 53155, 53156, 53157, 53158, 53159, 53160, 
    53161, 53162, 53163, 53164, 53165, 53166, 53167, 53168, 53169, 53170, 
    53171, 53172, 53173, 53174, 53175, 53176, 53177, 53178, 53179, 53180, 
    53181, 53182, 53183, 53184, 53185, 53186, 53187, 53188, 53189, 53190, 
    53191, 53192, 53193, 53194, 53195, 53196, 53197, 53198, 53199, 53200, 
    53201, 53202, 53203, 53204, 53205, 53206, 53207, 53208, 53209, 53210, 
    53211, 53212, 53213, 53214, 53215, 53216, 53217, 53218, 53219, 53220, 
    53221, 53222, 53223, 53224, 53225, 53226, 53227, 53228, 53229, 53230, 
    53231, 53232, 53233, 53234, 53235, 53236, 53237, 53238, 53239, 53240, 
    53241, 53242, 53243, 53244, 53245, 53246, 53247, 53248, 53249, 53250, 
    53251, 53252, 53253, 53254, 53255, 53256, 53257, 53258, 53259, 53260, 
    53261, 53262, 53263, 53264, 53265, 53266, 53267, 53268, 53269, 53270, 
    53271, 53272, 53273, 53274, 53275, 53276, 53277, 53278, 53279, 53280, 
    53281, 53282, 53283, 53284, 53285, 53286, 53287, 53288, 53289, 53290, 
    53291, 53292, 53293, 53294, 53295, 53296, 53297, 53298, 53299, 53300, 
    53301, 53302, 53303, 53304, 53305, 53306, 53307, 53308, 53309, 53310, 
    53311, 53312, 53313, 53314, 53315, 53316, 53317, 53318, 53319, 53320, 
    53321, 53322, 53323, 53324, 53325, 53326, 53327, 53328, 53329, 53330, 
    53331, 53332, 53333, 53334, 53335, 53336, 53337, 53338, 53339, 53340, 
    53341, 53342, 53343, 53344, 53345, 53346, 53347, 53348, 53349, 53350, 
    53351, 53352, 53353, 53354, 53355, 53356, 53357, 53358, 53359, 53360, 
    53361, 53362, 53363, 53364, 53365, 53366, 53367, 53368, 53369, 53370, 
    53371, 53372, 53373, 53374, 53375, 53376, 53377, 53378, 53379, 53380, 
    53381, 53382, 53383, 53384, 53385, 53386, 53387, 53388, 53389, 53390, 
    53391, 53392, 53393, 53394, 53395, 53396, 53397, 53398, 53399, 53400, 
    53401, 53402, 53403, 53404, 53405, 53406, 53407, 53408, 53409, 53410, 
    53411, 53412, 53413, 53414, 53415, 53416, 53417, 53418, 53419, 53420, 
    53421, 53422, 53423, 53424, 53425, 53426, 53427, 53428, 53429, 53430, 
    53431, 53432, 53433, 53434, 53435, 53436, 53437, 53438, 53439, 53440, 
    53441, 53442, 53443, 53444, 53445, 53446, 53447, 53448, 53449, 53450, 
    53451, 53452, 53453, 53454, 53455, 53456, 53457, 53458, 53459, 53460, 
    53461, 53462, 53463, 53464, 53465, 53466, 53467, 53468, 53469, 53470, 
    53471, 53472, 53473, 53474, 53475, 53476, 53477, 53478, 53479, 53480, 
    53481, 53482, 53483, 53484, 53485, 53486, 53487, 53488, 53489, 53490, 
    53491, 53492, 53493, 53494, 53495, 53496, 53497, 53498, 53499, 53500, 
    53501, 53502, 53503, 53504, 53505, 53506, 53507, 53508, 53509, 53510, 
    53511, 53512, 53513, 53514, 53515, 53516, 53517, 53518, 53519, 53520, 
    53521, 53522, 53523, 53524, 53525, 53526, 53527, 53528, 53529, 53530, 
    53531, 53532, 53533, 53534, 53535, 53536, 53537, 53538, 53539, 53540, 
    53541, 53542, 53543, 53544, 53545, 53546, 53547, 53548, 53549, 53550, 
    53551, 53552, 53553, 53554, 53555, 53556, 53557, 53558, 53559, 53560, 
    53561, 53562, 53563, 53564, 53565, 53566, 53567, 53568, 53569, 53570, 
    53571, 53572, 53573, 53574, 53575, 53576, 53577, 53578, 53579, 53580, 
    53581, 53582, 53583, 53584, 53585, 53586, 53587, 53588, 53589, 53590, 
    53591, 53592, 53593, 53594, 53595, 53596, 53597, 53598, 53599, 53600, 
    53601, 53602, 53603, 53604, 53605, 53606, 53607, 53608, 53609, 53610, 
    53611, 53612, 53613, 53614, 53615, 53616, 53617, 53618, 53619, 53620, 
    53621, 53622, 53623, 53624, 53625, 53626, 53627, 53628, 53629, 53630, 
    53631, 53632, 53633, 53634, 53635, 53636, 53637, 53638, 53639, 53640, 
    53641, 53642, 53643, 53644, 53645, 53646, 53647, 53648, 53649, 53650, 
    53651, 53652, 53653, 53654, 53655, 53656, 53657, 53658, 53659, 53660, 
    53661, 53662, 53663, 53664, 53665, 53666, 53667, 53668, 53669, 53670, 
    53671, 53672, 53673, 53674, 53675, 53676, 53677, 53678, 53679, 53680, 
    53681, 53682, 53683, 53684, 53685, 53686, 53687, 53688, 53689, 53690, 
    53691, 53692, 53693, 53694, 53695, 53696, 53697, 53698, 53699, 53700, 
    53701, 53702, 53703, 53704, 53705, 53706, 53707, 53708, 53709, 53710, 
    53711, 53712, 53713, 53714, 53715, 53716, 53717, 53718, 53719, 53720, 
    53721, 53722, 53723, 53724, 53725, 53726, 53727, 53728, 53729, 53730, 
    53731, 53732, 53733, 53734, 53735, 53736, 53737, 53738, 53739, 53740, 
    53741, 53742, 53743, 53744, 53745, 53746, 53747, 53748, 53749, 53750, 
    53751, 53752, 53753, 53754, 53755, 53756, 53757, 53758, 53759, 53760, 
    53761, 53762, 53763, 53764, 53765, 53766, 53767, 53768, 53769, 53770, 
    53771, 53772, 53773, 53774, 53775, 53776, 53777, 53778, 53779, 53780, 
    53781, 53782, 53783, 53784, 53785, 53786, 53787, 53788, 53789, 53790, 
    53791, 53792, 53793, 53794, 53795, 53796, 53797, 53798, 53799, 53800, 
    53801, 53802, 53803, 53804, 53805, 53806, 53807, 53808, 53809, 53810, 
    53811, 53812, 53813, 53814, 53815, 53816, 53817, 53818, 53819, 53820, 
    53821, 53822, 53823, 53824, 53825, 53826, 53827, 53828, 53829, 53830, 
    53831, 53832, 53833, 53834, 53835, 53836, 53837, 53838, 53839, 53840, 
    53841, 53842, 53843, 53844, 53845, 53846, 53847, 53848, 53849, 53850, 
    53851, 53852, 53853, 53854, 53855, 53856, 53857, 53858, 53859, 53860, 
    53861, 53862, 53863, 53864, 53865, 53866, 53867, 53868, 53869, 53870, 
    53871, 53872, 53873, 53874, 53875, 53876, 53877, 53878, 53879, 53880, 
    53881, 53882, 53883, 53884, 53885, 53886, 53887, 53888, 53889, 53890, 
    53891, 53892, 53893, 53894, 53895, 53896, 53897, 53898, 53899, 53900, 
    53901, 53902, 53903, 53904, 53905, 53906, 53907, 53908, 53909, 53910, 
    53911, 53912, 53913, 53914, 53915, 53916, 53917, 53918, 53919, 53920, 
    53921, 53922, 53923, 53924, 53925, 53926, 53927, 53928, 53929, 53930, 
    53931, 53932, 53933, 53934, 53935, 53936, 53937, 53938, 53939, 53940, 
    53941, 53942, 53943, 53944, 53945, 53946, 53947, 53948, 53949, 53950, 
    53951, 53952, 53953, 53954, 53955, 53956, 53957, 53958, 53959, 53960, 
    53961, 53962, 53963, 53964, 53965, 53966, 53967, 53968, 53969, 53970, 
    53971, 53972, 53973, 53974, 53975, 53976, 53977, 53978, 53979, 53980, 
    53981, 53982, 53983, 53984, 53985, 53986, 53987, 53988, 53989, 53990, 
    53991, 53992, 53993, 53994, 53995, 53996, 53997, 53998, 53999, 54000, 
    54001, 54002, 54003, 54004, 54005, 54006, 54007, 54008, 54009, 54010, 
    54011, 54012, 54013, 54014, 54015, 54016, 54017, 54018, 54019, 54020, 
    54021, 54022, 54023, 54024, 54025, 54026, 54027, 54028, 54029, 54030, 
    54031, 54032, 54033, 54034, 54035, 54036, 54037, 54038, 54039, 54040, 
    54041, 54042, 54043, 54044, 54045, 54046, 54047, 54048, 54049, 54050, 
    54051, 54052, 54053, 54054, 54055, 54056, 54057, 54058, 54059, 54060, 
    54061, 54062, 54063, 54064, 54065, 54066, 54067, 54068, 54069, 54070, 
    54071, 54072, 54073, 54074, 54075, 54076, 54077, 54078, 54079, 54080, 
    54081, 54082, 54083, 54084, 54085, 54086, 54087, 54088, 54089, 54090, 
    54091, 54092, 54093, 54094, 54095, 54096, 54097, 54098, 54099, 54100, 
    54101, 54102, 54103, 54104, 54105, 54106, 54107, 54108, 54109, 54110, 
    54111, 54112, 54113, 54114, 54115, 54116, 54117, 54118, 54119, 54120, 
    54121, 54122, 54123, 54124, 54125, 54126, 54127, 54128, 54129, 54130, 
    54131, 54132, 54133, 54134, 54135, 54136, 54137, 54138, 54139, 54140, 
    54141, 54142, 54143, 54144, 54145, 54146, 54147, 54148, 54149, 54150, 
    54151, 54152, 54153, 54154, 54155, 54156, 54157, 54158, 54159, 54160, 
    54161, 54162, 54163, 54164, 54165, 54166, 54167, 54168, 54169, 54170, 
    54171, 54172, 54173, 54174, 54175, 54176, 54177, 54178, 54179, 54180, 
    54181, 54182, 54183, 54184, 54185, 54186, 54187, 54188, 54189, 54190, 
    54191, 54192, 54193, 54194, 54195, 54196, 54197, 54198, 54199, 54200, 
    54201, 54202, 54203, 54204, 54205, 54206, 54207, 54208, 54209, 54210, 
    54211, 54212, 54213, 54214, 54215, 54216, 54217, 54218, 54219, 54220, 
    54221, 54222, 54223, 54224, 54225, 54226, 54227, 54228, 54229, 54230, 
    54231, 54232, 54233, 54234, 54235, 54236, 54237, 54238, 54239, 54240, 
    54241, 54242, 54243, 54244, 54245, 54246, 54247, 54248, 54249, 54250, 
    54251, 54252, 54253, 54254, 54255, 54256, 54257, 54258, 54259, 54260, 
    54261, 54262, 54263, 54264, 54265, 54266, 54267, 54268, 54269, 54270, 
    54271, 54272, 54273, 54274, 54275, 54276, 54277, 54278, 54279, 54280, 
    54281, 54282, 54283, 54284, 54285, 54286, 54287, 54288, 54289, 54290, 
    54291, 54292, 54293, 54294, 54295, 54296, 54297, 54298, 54299, 54300, 
    54301, 54302, 54303, 54304, 54305, 54306, 54307, 54308, 54309, 54310, 
    54311, 54312, 54313, 54314, 54315, 54316, 54317, 54318, 54319, 54320, 
    54321, 54322, 54323, 54324, 54325, 54326, 54327, 54328, 54329, 54330, 
    54331, 54332, 54333, 54334, 54335, 54336, 54337, 54338, 54339, 54340, 
    54341, 54342, 54343, 54344, 54345, 54346, 54347, 54348, 54349, 54350, 
    54351, 54352, 54353, 54354, 54355, 54356, 54357, 54358, 54359, 54360, 
    54361, 54362, 54363, 54364, 54365, 54366, 54367, 54368, 54369, 54370, 
    54371, 54372, 54373, 54374, 54375, 54376, 54377, 54378, 54379, 54380, 
    54381, 54382, 54383, 54384, 54385, 54386, 54387, 54388, 54389, 54390, 
    54391, 54392, 54393, 54394, 54395, 54396, 54397, 54398, 54399, 54400, 
    54401, 54402, 54403, 54404, 54405, 54406, 54407, 54408, 54409, 54410, 
    54411, 54412, 54413, 54414, 54415, 54416, 54417, 54418, 54419, 54420, 
    54421, 54422, 54423, 54424, 54425, 54426, 54427, 54428, 54429, 54430, 
    54431, 54432, 54433, 54434, 54435, 54436, 54437, 54438, 54439, 54440, 
    54441, 54442, 54443, 54444, 54445, 54446, 54447, 54448, 54449, 54450, 
    54451, 54452, 54453, 54454, 54455, 54456, 54457, 54458, 54459, 54460, 
    54461, 54462, 54463, 54464, 54465, 54466, 54467, 54468, 54469, 54470, 
    54471, 54472, 54473, 54474, 54475, 54476, 54477, 54478, 54479, 54480, 
    54481, 54482, 54483, 54484, 54485, 54486, 54487, 54488, 54489, 54490, 
    54491, 54492, 54493, 54494, 54495, 54496, 54497, 54498, 54499, 54500, 
    54501, 54502, 54503, 54504, 54505, 54506, 54507, 54508, 54509, 54510, 
    54511, 54512, 54513, 54514, 54515, 54516, 54517, 54518, 54519, 54520, 
    54521, 54522, 54523, 54524, 54525, 54526, 54527, 54528, 54529, 54530, 
    54531, 54532, 54533, 54534, 54535, 54536, 54537, 54538, 54539, 54540, 
    54541, 54542, 54543, 54544, 54545, 54546, 54547, 54548, 54549, 54550, 
    54551, 54552, 54553, 54554, 54555, 54556, 54557, 54558, 54559, 54560, 
    54561, 54562, 54563, 54564, 54565, 54566, 54567, 54568, 54569, 54570, 
    54571, 54572, 54573, 54574, 54575, 54576, 54577, 54578, 54579, 54580, 
    54581, 54582, 54583, 54584, 54585, 54586, 54587, 54588, 54589, 54590, 
    54591, 54592, 54593, 54594, 54595, 54596, 54597, 54598, 54599, 54600, 
    54601, 54602, 54603, 54604, 54605, 54606, 54607, 54608, 54609, 54610, 
    54611, 54612, 54613, 54614, 54615, 54616, 54617, 54618, 54619, 54620, 
    54621, 54622, 54623, 54624, 54625, 54626, 54627, 54628, 54629, 54630, 
    54631, 54632, 54633, 54634, 54635, 54636, 54637, 54638, 54639, 54640, 
    54641, 54642, 54643, 54644, 54645, 54646, 54647, 54648, 54649, 54650, 
    54651, 54652, 54653, 54654, 54655, 54656, 54657, 54658, 54659, 54660, 
    54661, 54662, 54663, 54664, 54665, 54666, 54667, 54668, 54669, 54670, 
    54671, 54672, 54673, 54674, 54675, 54676, 54677, 54678, 54679, 54680, 
    54681, 54682, 54683, 54684, 54685, 54686, 54687, 54688, 54689, 54690, 
    54691, 54692, 54693, 54694, 54695, 54696, 54697, 54698, 54699, 54700, 
    54701, 54702, 54703, 54704, 54705, 54706, 54707, 54708, 54709, 54710, 
    54711, 54712, 54713, 54714, 54715, 54716, 54717, 54718, 54719, 54720, 
    54721, 54722, 54723, 54724, 54725, 54726, 54727, 54728, 54729, 54730, 
    54731, 54732, 54733, 54734, 54735, 54736, 54737, 54738, 54739, 54740, 
    54741, 54742, 54743, 54744, 54745, 54746, 54747, 54748, 54749, 54750, 
    54751, 54752, 54753, 54754, 54755, 54756, 54757, 54758, 54759, 54760, 
    54761, 54762, 54763, 54764, 54765, 54766, 54767, 54768, 54769, 54770, 
    54771, 54772, 54773, 54774, 54775, 54776, 54777, 54778, 54779, 54780, 
    54781, 54782, 54783, 54784, 54785, 54786, 54787, 54788, 54789, 54790, 
    54791, 54792, 54793, 54794, 54795, 54796, 54797, 54798, 54799, 54800, 
    54801, 54802, 54803, 54804, 54805, 54806, 54807, 54808, 54809, 54810, 
    54811, 54812, 54813, 54814, 54815, 54816, 54817, 54818, 54819, 54820, 
    54821, 54822, 54823, 54824, 54825, 54826, 54827, 54828, 54829, 54830, 
    54831, 54832, 54833, 54834, 54835, 54836, 54837, 54838, 54839, 54840, 
    54841, 54842, 54843, 54844, 54845, 54846, 54847, 54848, 54849, 54850, 
    54851, 54852, 54853, 54854, 54855, 54856, 54857, 54858, 54859, 54860, 
    54861, 54862, 54863, 54864, 54865, 54866, 54867, 54868, 54869, 54870, 
    54871, 54872, 54873, 54874, 54875, 54876, 54877, 54878, 54879, 54880, 
    54881, 54882, 54883, 54884, 54885, 54886, 54887, 54888, 54889, 54890, 
    54891, 54892, 54893, 54894, 54895, 54896, 54897, 54898, 54899, 54900, 
    54901, 54902, 54903, 54904, 54905, 54906, 54907, 54908, 54909, 54910, 
    54911, 54912, 54913, 54914, 54915, 54916, 54917, 54918, 54919, 54920, 
    54921, 54922, 54923, 54924, 54925, 54926, 54927, 54928, 54929, 54930, 
    54931, 54932, 54933, 54934, 54935, 54936, 54937, 54938, 54939, 54940, 
    54941, 54942, 54943, 54944, 54945, 54946, 54947, 54948, 54949, 54950, 
    54951, 54952, 54953, 54954, 54955, 54956, 54957, 54958, 54959, 54960, 
    54961, 54962, 54963, 54964, 54965, 54966, 54967, 54968, 54969, 54970, 
    54971, 54972, 54973, 54974, 54975, 54976, 54977, 54978, 54979, 54980, 
    54981, 54982, 54983, 54984, 54985, 54986, 54987, 54988, 54989, 54990, 
    54991, 54992, 54993, 54994, 54995, 54996, 54997, 54998, 54999, 55000, 
    55001, 55002, 55003, 55004, 55005, 55006, 55007, 55008, 55009, 55010, 
    55011, 55012, 55013, 55014, 55015, 55016, 55017, 55018, 55019, 55020, 
    55021, 55022, 55023, 55024, 55025, 55026, 55027, 55028, 55029, 55030, 
    55031, 55032, 55033, 55034, 55035, 55036, 55037, 55038, 55039, 55040, 
    55041, 55042, 55043, 55044, 55045, 55046, 55047, 55048, 55049, 55050, 
    55051, 55052, 55053, 55054, 55055, 55056, 55057, 55058, 55059, 55060, 
    55061, 55062, 55063, 55064, 55065, 55066, 55067, 55068, 55069, 55070, 
    55071, 55072, 55073, 55074, 55075, 55076, 55077, 55078, 55079, 55080, 
    55081, 55082, 55083, 55084, 55085, 55086, 55087, 55088, 55089, 55090, 
    55091, 55092, 55093, 55094, 55095, 55096, 55097, 55098, 55099, 55100, 
    55101, 55102, 55103, 55104, 55105, 55106, 55107, 55108, 55109, 55110, 
    55111, 55112, 55113, 55114, 55115, 55116, 55117, 55118, 55119, 55120, 
    55121, 55122, 55123, 55124, 55125, 55126, 55127, 55128, 55129, 55130, 
    55131, 55132, 55133, 55134, 55135, 55136, 55137, 55138, 55139, 55140, 
    55141, 55142, 55143, 55144, 55145, 55146, 55147, 55148, 55149, 55150, 
    55151, 55152, 55153, 55154, 55155, 55156, 55157, 55158, 55159, 55160, 
    55161, 55162, 55163, 55164, 55165, 55166, 55167, 55168, 55169, 55170, 
    55171, 55172, 55173, 55174, 55175, 55176, 55177, 55178, 55179, 55180, 
    55181, 55182, 55183, 55184, 55185, 55186, 55187, 55188, 55189, 55190, 
    55191, 55192, 55193, 55194, 55195, 55196, 55197, 55198, 55199, 55200, 
    55201, 55202, 55203, 55204, 55205, 55206, 55207, 55208, 55209, 55210, 
    55211, 55212, 55213, 55214, 55215, 55216, 55217, 55218, 55219, 55220, 
    55221, 55222, 55223, 55224, 55225, 55226, 55227, 55228, 55229, 55230, 
    55231, 55232, 55233, 55234, 55235, 55236, 55237, 55238, 55239, 55240, 
    55241, 55242, 55243, 55244, 55245, 55246, 55247, 55248, 55249, 55250, 
    55251, 55252, 55253, 55254, 55255, 55256, 55257, 55258, 55259, 55260, 
    55261, 55262, 55263, 55264, 55265, 55266, 55267, 55268, 55269, 55270, 
    55271, 55272, 55273, 55274, 55275, 55276, 55277, 55278, 55279, 55280, 
    55281, 55282, 55283, 55284, 55285, 55286, 55287, 55288, 55289, 55290, 
    55291, 55292, 55293, 55294, 55295, 55296, 55297, 55298, 55299, 55300, 
    55301, 55302, 55303, 55304, 55305, 55306, 55307, 55308, 55309, 55310, 
    55311, 55312, 55313, 55314, 55315, 55316, 55317, 55318, 55319, 55320, 
    55321, 55322, 55323, 55324, 55325, 55326, 55327, 55328, 55329, 55330, 
    55331, 55332, 55333, 55334, 55335, 55336, 55337, 55338, 55339, 55340, 
    55341, 55342, 55343, 55344, 55345, 55346, 55347, 55348, 55349, 55350, 
    55351, 55352, 55353, 55354, 55355, 55356, 55357, 55358, 55359, 55360, 
    55361, 55362, 55363, 55364, 55365, 55366, 55367, 55368, 55369, 55370, 
    55371, 55372, 55373, 55374, 55375, 55376, 55377, 55378, 55379, 55380, 
    55381, 55382, 55383, 55384, 55385, 55386, 55387, 55388, 55389, 55390, 
    55391, 55392, 55393, 55394, 55395, 55396, 55397, 55398, 55399, 55400, 
    55401, 55402, 55403, 55404, 55405, 55406, 55407, 55408, 55409, 55410, 
    55411, 55412, 55413, 55414, 55415, 55416, 55417, 55418, 55419, 55420, 
    55421, 55422, 55423, 55424, 55425, 55426, 55427, 55428, 55429, 55430, 
    55431, 55432, 55433, 55434, 55435, 55436, 55437, 55438, 55439, 55440, 
    55441, 55442, 55443, 55444, 55445, 55446, 55447, 55448, 55449, 55450, 
    55451, 55452, 55453, 55454, 55455, 55456, 55457, 55458, 55459, 55460, 
    55461, 55462, 55463, 55464, 55465, 55466, 55467, 55468, 55469, 55470, 
    55471, 55472, 55473, 55474, 55475, 55476, 55477, 55478, 55479, 55480, 
    55481, 55482, 55483, 55484, 55485, 55486, 55487, 55488, 55489, 55490, 
    55491, 55492, 55493, 55494, 55495, 55496, 55497, 55498, 55499, 55500, 
    55501, 55502, 55503, 55504, 55505, 55506, 55507, 55508, 55509, 55510, 
    55511, 55512, 55513, 55514, 55515, 55516, 55517, 55518, 55519, 55520, 
    55521, 55522, 55523, 55524, 55525, 55526, 55527, 55528, 55529, 55530, 
    55531, 55532, 55533, 55534, 55535, 55536, 55537, 55538, 55539, 55540, 
    55541, 55542, 55543, 55544, 55545, 55546, 55547, 55548, 55549, 55550, 
    55551, 55552, 55553, 55554, 55555, 55556, 55557, 55558, 55559, 55560, 
    55561, 55562, 55563, 55564, 55565, 55566, 55567, 55568, 55569, 55570, 
    55571, 55572, 55573, 55574, 55575, 55576, 55577, 55578, 55579, 55580, 
    55581, 55582, 55583, 55584, 55585, 55586, 55587, 55588, 55589, 55590, 
    55591, 55592, 55593, 55594, 55595, 55596, 55597, 55598, 55599, 55600, 
    55601, 55602, 55603, 55604, 55605, 55606, 55607, 55608, 55609, 55610, 
    55611, 55612, 55613, 55614, 55615, 55616, 55617, 55618, 55619, 55620, 
    55621, 55622, 55623, 55624, 55625, 55626, 55627, 55628, 55629, 55630, 
    55631, 55632, 55633, 55634, 55635, 55636, 55637, 55638, 55639, 55640, 
    55641, 55642, 55643, 55644, 55645, 55646, 55647, 55648, 55649, 55650, 
    55651, 55652, 55653, 55654, 55655, 55656, 55657, 55658, 55659, 55660, 
    55661, 55662, 55663, 55664, 55665, 55666, 55667, 55668, 55669, 55670, 
    55671, 55672, 55673, 55674, 55675, 55676, 55677, 55678, 55679, 55680, 
    55681, 55682, 55683, 55684, 55685, 55686, 55687, 55688, 55689, 55690, 
    55691, 55692, 55693, 55694, 55695, 55696, 55697, 55698, 55699, 55700, 
    55701, 55702, 55703, 55704, 55705, 55706, 55707, 55708, 55709, 55710, 
    55711, 55712, 55713, 55714, 55715, 55716, 55717, 55718, 55719, 55720, 
    55721, 55722, 55723, 55724, 55725, 55726, 55727, 55728, 55729, 55730, 
    55731, 55732, 55733, 55734, 55735, 55736, 55737, 55738, 55739, 55740, 
    55741, 55742, 55743, 55744, 55745, 55746, 55747, 55748, 55749, 55750, 
    55751, 55752, 55753, 55754, 55755, 55756, 55757, 55758, 55759, 55760, 
    55761, 55762, 55763, 55764, 55765, 55766, 55767, 55768, 55769, 55770, 
    55771, 55772, 55773, 55774, 55775, 55776, 55777, 55778, 55779, 55780, 
    55781, 55782, 55783, 55784, 55785, 55786, 55787, 55788, 55789, 55790, 
    55791, 55792, 55793, 55794, 55795, 55796, 55797, 55798, 55799, 55800, 
    55801, 55802, 55803, 55804, 55805, 55806, 55807, 55808, 55809, 55810, 
    55811, 55812, 55813, 55814, 55815, 55816, 55817, 55818, 55819, 55820, 
    55821, 55822, 55823, 55824, 55825, 55826, 55827, 55828, 55829, 55830, 
    55831, 55832, 55833, 55834, 55835, 55836, 55837, 55838, 55839, 55840, 
    55841, 55842, 55843, 55844, 55845, 55846, 55847, 55848, 55849, 55850, 
    55851, 55852, 55853, 55854, 55855, 55856, 55857, 55858, 55859, 55860, 
    55861, 55862, 55863, 55864, 55865, 55866, 55867, 55868, 55869, 55870, 
    55871, 55872, 55873, 55874, 55875, 55876, 55877, 55878, 55879, 55880, 
    55881, 55882, 55883, 55884, 55885, 55886, 55887, 55888, 55889, 55890, 
    55891, 55892, 55893, 55894, 55895, 55896, 55897, 55898, 55899, 55900, 
    55901, 55902, 55903, 55904, 55905, 55906, 55907, 55908, 55909, 55910, 
    55911, 55912, 55913, 55914, 55915, 55916, 55917, 55918, 55919, 55920, 
    55921, 55922, 55923, 55924, 55925, 55926, 55927, 55928, 55929, 55930, 
    55931, 55932, 55933, 55934, 55935, 55936, 55937, 55938, 55939, 55940, 
    55941, 55942, 55943, 55944, 55945, 55946, 55947, 55948, 55949, 55950, 
    55951, 55952, 55953, 55954, 55955, 55956, 55957, 55958, 55959, 55960, 
    55961, 55962, 55963, 55964, 55965, 55966, 55967, 55968, 55969, 55970, 
    55971, 55972, 55973, 55974, 55975, 55976, 55977, 55978, 55979, 55980, 
    55981, 55982, 55983, 55984, 55985, 55986, 55987, 55988, 55989, 55990, 
    55991, 55992, 55993, 55994, 55995, 55996, 55997, 55998, 55999, 56000, 
    56001, 56002, 56003, 56004, 56005, 56006, 56007, 56008, 56009, 56010, 
    56011, 56012, 56013, 56014, 56015, 56016, 56017, 56018, 56019, 56020, 
    56021, 56022, 56023, 56024, 56025, 56026, 56027, 56028, 56029, 56030, 
    56031, 56032, 56033, 56034, 56035, 56036, 56037, 56038, 56039, 56040, 
    56041, 56042, 56043, 56044, 56045, 56046, 56047, 56048, 56049, 56050, 
    56051, 56052, 56053, 56054, 56055, 56056, 56057, 56058, 56059, 56060, 
    56061, 56062, 56063, 56064, 56065, 56066, 56067, 56068, 56069, 56070, 
    56071, 56072, 56073, 56074, 56075, 56076, 56077, 56078, 56079, 56080, 
    56081, 56082, 56083, 56084, 56085, 56086, 56087, 56088, 56089, 56090, 
    56091, 56092, 56093, 56094, 56095, 56096, 56097, 56098, 56099, 56100, 
    56101, 56102, 56103, 56104, 56105, 56106, 56107, 56108, 56109, 56110, 
    56111, 56112, 56113, 56114, 56115, 56116, 56117, 56118, 56119, 56120, 
    56121, 56122, 56123, 56124, 56125, 56126, 56127, 56128, 56129, 56130, 
    56131, 56132, 56133, 56134, 56135, 56136, 56137, 56138, 56139, 56140, 
    56141, 56142, 56143, 56144, 56145, 56146, 56147, 56148, 56149, 56150, 
    56151, 56152, 56153, 56154, 56155, 56156, 56157, 56158, 56159, 56160, 
    56161, 56162, 56163, 56164, 56165, 56166, 56167, 56168, 56169, 56170, 
    56171, 56172, 56173, 56174, 56175, 56176, 56177, 56178, 56179, 56180, 
    56181, 56182, 56183, 56184, 56185, 56186, 56187, 56188, 56189, 56190, 
    56191, 56192, 56193, 56194, 56195, 56196, 56197, 56198, 56199, 56200, 
    56201, 56202, 56203, 56204, 56205, 56206, 56207, 56208, 56209, 56210, 
    56211, 56212, 56213, 56214, 56215, 56216, 56217, 56218, 56219, 56220, 
    56221, 56222, 56223, 56224, 56225, 56226, 56227, 56228, 56229, 56230, 
    56231, 56232, 56233, 56234, 56235, 56236, 56237, 56238, 56239, 56240, 
    56241, 56242, 56243, 56244, 56245, 56246, 56247, 56248, 56249, 56250, 
    56251, 56252, 56253, 56254, 56255, 56256, 56257, 56258, 56259, 56260, 
    56261, 56262, 56263, 56264, 56265, 56266, 56267, 56268, 56269, 56270, 
    56271, 56272, 56273, 56274, 56275, 56276, 56277, 56278, 56279, 56280, 
    56281, 56282, 56283, 56284, 56285, 56286, 56287, 56288, 56289, 56290, 
    56291, 56292, 56293, 56294, 56295, 56296, 56297, 56298, 56299, 56300, 
    56301, 56302, 56303, 56304, 56305, 56306, 56307, 56308, 56309, 56310, 
    56311, 56312, 56313, 56314, 56315, 56316, 56317, 56318, 56319, 56320, 
    56321, 56322, 56323, 56324, 56325, 56326, 56327, 56328, 56329, 56330, 
    56331, 56332, 56333, 56334, 56335, 56336, 56337, 56338, 56339, 56340, 
    56341, 56342, 56343, 56344, 56345, 56346, 56347, 56348, 56349, 56350, 
    56351, 56352, 56353, 56354, 56355, 56356, 56357, 56358, 56359, 56360, 
    56361, 56362, 56363, 56364, 56365, 56366, 56367, 56368, 56369, 56370, 
    56371, 56372, 56373, 56374, 56375, 56376, 56377, 56378, 56379, 56380, 
    56381, 56382, 56383, 56384, 56385, 56386, 56387, 56388, 56389, 56390, 
    56391, 56392, 56393, 56394, 56395, 56396, 56397, 56398, 56399, 56400, 
    56401, 56402, 56403, 56404, 56405, 56406, 56407, 56408, 56409, 56410, 
    56411, 56412, 56413, 56414, 56415, 56416, 56417, 56418, 56419, 56420, 
    56421, 56422, 56423, 56424, 56425, 56426, 56427, 56428, 56429, 56430, 
    56431, 56432, 56433, 56434, 56435, 56436, 56437, 56438, 56439, 56440, 
    56441, 56442, 56443, 56444, 56445, 56446, 56447, 56448, 56449, 56450, 
    56451, 56452, 56453, 56454, 56455, 56456, 56457, 56458, 56459, 56460, 
    56461, 56462, 56463, 56464, 56465, 56466, 56467, 56468, 56469, 56470, 
    56471, 56472, 56473, 56474, 56475, 56476, 56477, 56478, 56479, 56480, 
    56481, 56482, 56483, 56484, 56485, 56486, 56487, 56488, 56489, 56490, 
    56491, 56492, 56493, 56494, 56495, 56496, 56497, 56498, 56499, 56500, 
    56501, 56502, 56503, 56504, 56505, 56506, 56507, 56508, 56509, 56510, 
    56511, 56512, 56513, 56514, 56515, 56516, 56517, 56518, 56519, 56520, 
    56521, 56522, 56523, 56524, 56525, 56526, 56527, 56528, 56529, 56530, 
    56531, 56532, 56533, 56534, 56535, 56536, 56537, 56538, 56539, 56540, 
    56541, 56542, 56543, 56544, 56545, 56546, 56547, 56548, 56549, 56550, 
    56551, 56552, 56553, 56554, 56555, 56556, 56557, 56558, 56559, 56560, 
    56561, 56562, 56563, 56564, 56565, 56566, 56567, 56568, 56569, 56570, 
    56571, 56572, 56573, 56574, 56575, 56576, 56577, 56578, 56579, 56580, 
    56581, 56582, 56583, 56584, 56585, 56586, 56587, 56588, 56589, 56590, 
    56591, 56592, 56593, 56594, 56595, 56596, 56597, 56598, 56599, 56600, 
    56601, 56602, 56603, 56604, 56605, 56606, 56607, 56608, 56609, 56610, 
    56611, 56612, 56613, 56614, 56615, 56616, 56617, 56618, 56619, 56620, 
    56621, 56622, 56623, 56624, 56625, 56626, 56627, 56628, 56629, 56630, 
    56631, 56632, 56633, 56634, 56635, 56636, 56637, 56638, 56639, 56640, 
    56641, 56642, 56643, 56644, 56645, 56646, 56647, 56648, 56649, 56650, 
    56651, 56652, 56653, 56654, 56655, 56656, 56657, 56658, 56659, 56660, 
    56661, 56662, 56663, 56664, 56665, 56666, 56667, 56668, 56669, 56670, 
    56671, 56672, 56673, 56674, 56675, 56676, 56677, 56678, 56679, 56680, 
    56681, 56682, 56683, 56684, 56685, 56686, 56687, 56688, 56689, 56690, 
    56691, 56692, 56693, 56694, 56695, 56696, 56697, 56698, 56699, 56700, 
    56701, 56702, 56703, 56704, 56705, 56706, 56707, 56708, 56709, 56710, 
    56711, 56712, 56713, 56714, 56715, 56716, 56717, 56718, 56719, 56720, 
    56721, 56722, 56723, 56724, 56725, 56726, 56727, 56728, 56729, 56730, 
    56731, 56732, 56733, 56734, 56735, 56736, 56737, 56738, 56739, 56740, 
    56741, 56742, 56743, 56744, 56745, 56746, 56747, 56748, 56749, 56750, 
    56751, 56752, 56753, 56754, 56755, 56756, 56757, 56758, 56759, 56760, 
    56761, 56762, 56763, 56764, 56765, 56766, 56767, 56768, 56769, 56770, 
    56771, 56772, 56773, 56774, 56775, 56776, 56777, 56778, 56779, 56780, 
    56781, 56782, 56783, 56784, 56785, 56786, 56787, 56788, 56789, 56790, 
    56791, 56792, 56793, 56794, 56795, 56796, 56797, 56798, 56799, 56800, 
    56801, 56802, 56803, 56804, 56805, 56806, 56807, 56808, 56809, 56810, 
    56811, 56812, 56813, 56814, 56815, 56816, 56817, 56818, 56819, 56820, 
    56821, 56822, 56823, 56824, 56825, 56826, 56827, 56828, 56829, 56830, 
    56831, 56832, 56833, 56834, 56835, 56836, 56837, 56838, 56839, 56840, 
    56841, 56842, 56843, 56844, 56845, 56846, 56847, 56848, 56849, 56850, 
    56851, 56852, 56853, 56854, 56855, 56856, 56857, 56858, 56859, 56860, 
    56861, 56862, 56863, 56864, 56865, 56866, 56867, 56868, 56869, 56870, 
    56871, 56872, 56873, 56874, 56875, 56876, 56877, 56878, 56879, 56880, 
    56881, 56882, 56883, 56884, 56885, 56886, 56887, 56888, 56889, 56890, 
    56891, 56892, 56893, 56894, 56895, 56896, 56897, 56898, 56899, 56900, 
    56901, 56902, 56903, 56904, 56905, 56906, 56907, 56908, 56909, 56910, 
    56911, 56912, 56913, 56914, 56915, 56916, 56917, 56918, 56919, 56920, 
    56921, 56922, 56923, 56924, 56925, 56926, 56927, 56928, 56929, 56930, 
    56931, 56932, 56933, 56934, 56935, 56936, 56937, 56938, 56939, 56940, 
    56941, 56942, 56943, 56944, 56945, 56946, 56947, 56948, 56949, 56950, 
    56951, 56952, 56953, 56954, 56955, 56956, 56957, 56958, 56959, 56960, 
    56961, 56962, 56963, 56964, 56965, 56966, 56967, 56968, 56969, 56970, 
    56971, 56972, 56973, 56974, 56975, 56976, 56977, 56978, 56979, 56980, 
    56981, 56982, 56983, 56984, 56985, 56986, 56987, 56988, 56989, 56990, 
    56991, 56992, 56993, 56994, 56995, 56996, 56997, 56998, 56999, 57000, 
    57001, 57002, 57003, 57004, 57005, 57006, 57007, 57008, 57009, 57010, 
    57011, 57012, 57013, 57014, 57015, 57016, 57017, 57018, 57019, 57020, 
    57021, 57022, 57023, 57024, 57025, 57026, 57027, 57028, 57029, 57030, 
    57031, 57032, 57033, 57034, 57035, 57036, 57037, 57038, 57039, 57040, 
    57041, 57042, 57043, 57044, 57045, 57046, 57047, 57048, 57049, 57050, 
    57051, 57052, 57053, 57054, 57055, 57056, 57057, 57058, 57059, 57060, 
    57061, 57062, 57063, 57064, 57065, 57066, 57067, 57068, 57069, 57070, 
    57071, 57072, 57073, 57074, 57075, 57076, 57077, 57078, 57079, 57080, 
    57081, 57082, 57083, 57084, 57085, 57086, 57087, 57088, 57089, 57090, 
    57091, 57092, 57093, 57094, 57095, 57096, 57097, 57098, 57099, 57100, 
    57101, 57102, 57103, 57104, 57105, 57106, 57107, 57108, 57109, 57110, 
    57111, 57112, 57113, 57114, 57115, 57116, 57117, 57118, 57119, 57120, 
    57121, 57122, 57123, 57124, 57125, 57126, 57127, 57128, 57129, 57130, 
    57131, 57132, 57133, 57134, 57135, 57136, 57137, 57138, 57139, 57140, 
    57141, 57142, 57143, 57144, 57145, 57146, 57147, 57148, 57149, 57150, 
    57151, 57152, 57153, 57154, 57155, 57156, 57157, 57158, 57159, 57160, 
    57161, 57162, 57163, 57164, 57165, 57166, 57167, 57168, 57169, 57170, 
    57171, 57172, 57173, 57174, 57175, 57176, 57177, 57178, 57179, 57180, 
    57181, 57182, 57183, 57184, 57185, 57186, 57187, 57188, 57189, 57190, 
    57191, 57192, 57193, 57194, 57195, 57196, 57197, 57198, 57199, 57200, 
    57201, 57202, 57203, 57204, 57205, 57206, 57207, 57208, 57209, 57210, 
    57211, 57212, 57213, 57214, 57215, 57216, 57217, 57218, 57219, 57220, 
    57221, 57222, 57223, 57224, 57225, 57226, 57227, 57228, 57229, 57230, 
    57231, 57232, 57233, 57234, 57235, 57236, 57237, 57238, 57239, 57240, 
    57241, 57242, 57243, 57244, 57245, 57246, 57247, 57248, 57249, 57250, 
    57251, 57252, 57253, 57254, 57255, 57256, 57257, 57258, 57259, 57260, 
    57261, 57262, 57263, 57264, 57265, 57266, 57267, 57268, 57269, 57270, 
    57271, 57272, 57273, 57274, 57275, 57276, 57277, 57278, 57279, 57280, 
    57281, 57282, 57283, 57284, 57285, 57286, 57287, 57288, 57289, 57290, 
    57291, 57292, 57293, 57294, 57295, 57296, 57297, 57298, 57299, 57300, 
    57301, 57302, 57303, 57304, 57305, 57306, 57307, 57308, 57309, 57310, 
    57311, 57312, 57313, 57314, 57315, 57316, 57317, 57318, 57319, 57320, 
    57321, 57322, 57323, 57324, 57325, 57326, 57327, 57328, 57329, 57330, 
    57331, 57332, 57333, 57334, 57335, 57336, 57337, 57338, 57339, 57340, 
    57341, 57342, 57343, 57344, 57345, 57346, 57347, 57348, 57349, 57350, 
    57351, 57352, 57353, 57354, 57355, 57356, 57357, 57358, 57359, 57360, 
    57361, 57362, 57363, 57364, 57365, 57366, 57367, 57368, 57369, 57370, 
    57371, 57372, 57373, 57374, 57375, 57376, 57377, 57378, 57379, 57380, 
    57381, 57382, 57383, 57384, 57385, 57386, 57387, 57388, 57389, 57390, 
    57391, 57392, 57393, 57394, 57395, 57396, 57397, 57398, 57399, 57400, 
    57401, 57402, 57403, 57404, 57405, 57406, 57407, 57408, 57409, 57410, 
    57411, 57412, 57413, 57414, 57415, 57416, 57417, 57418, 57419, 57420, 
    57421, 57422, 57423, 57424, 57425, 57426, 57427, 57428, 57429, 57430, 
    57431, 57432, 57433, 57434, 57435, 57436, 57437, 57438, 57439, 57440, 
    57441, 57442, 57443, 57444, 57445, 57446, 57447, 57448, 57449, 57450, 
    57451, 57452, 57453, 57454, 57455, 57456, 57457, 57458, 57459, 57460, 
    57461, 57462, 57463, 57464, 57465, 57466, 57467, 57468, 57469, 57470, 
    57471, 57472, 57473, 57474, 57475, 57476, 57477, 57478, 57479, 57480, 
    57481, 57482, 57483, 57484, 57485, 57486, 57487, 57488, 57489, 57490, 
    57491, 57492, 57493, 57494, 57495, 57496, 57497, 57498, 57499, 57500, 
    57501, 57502, 57503, 57504, 57505, 57506, 57507, 57508, 57509, 57510, 
    57511, 57512, 57513, 57514, 57515, 57516, 57517, 57518, 57519, 57520, 
    57521, 57522, 57523, 57524, 57525, 57526, 57527, 57528, 57529, 57530, 
    57531, 57532, 57533, 57534, 57535, 57536, 57537, 57538, 57539, 57540, 
    57541, 57542, 57543, 57544, 57545, 57546, 57547, 57548, 57549, 57550, 
    57551, 57552, 57553, 57554, 57555, 57556, 57557, 57558, 57559, 57560, 
    57561, 57562, 57563, 57564, 57565, 57566, 57567, 57568, 57569, 57570, 
    57571, 57572, 57573, 57574, 57575, 57576, 57577, 57578, 57579, 57580, 
    57581, 57582, 57583, 57584, 57585, 57586, 57587, 57588, 57589, 57590, 
    57591, 57592, 57593, 57594, 57595, 57596, 57597, 57598, 57599, 57600, 
    57601, 57602, 57603, 57604, 57605, 57606, 57607, 57608, 57609, 57610, 
    57611, 57612, 57613, 57614, 57615, 57616, 57617, 57618, 57619, 57620, 
    57621, 57622, 57623, 57624, 57625, 57626, 57627, 57628, 57629, 57630, 
    57631, 57632, 57633, 57634, 57635, 57636, 57637, 57638, 57639, 57640, 
    57641, 57642, 57643, 57644, 57645, 57646, 57647, 57648, 57649, 57650, 
    57651, 57652, 57653, 57654, 57655, 57656, 57657, 57658, 57659, 57660, 
    57661, 57662, 57663, 57664, 57665, 57666, 57667, 57668, 57669, 57670, 
    57671, 57672, 57673, 57674, 57675, 57676, 57677, 57678, 57679, 57680, 
    57681, 57682, 57683, 57684, 57685, 57686, 57687, 57688, 57689, 57690, 
    57691, 57692, 57693, 57694, 57695, 57696, 57697, 57698, 57699, 57700, 
    57701, 57702, 57703, 57704, 57705, 57706, 57707, 57708, 57709, 57710, 
    57711, 57712, 57713, 57714, 57715, 57716, 57717, 57718, 57719, 57720, 
    57721, 57722, 57723, 57724, 57725, 57726, 57727, 57728, 57729, 57730, 
    57731, 57732, 57733, 57734, 57735, 57736, 57737, 57738, 57739, 57740, 
    57741, 57742, 57743, 57744, 57745, 57746, 57747, 57748, 57749, 57750, 
    57751, 57752, 57753, 57754, 57755, 57756, 57757, 57758, 57759, 57760, 
    57761, 57762, 57763, 57764, 57765, 57766, 57767, 57768, 57769, 57770, 
    57771, 57772, 57773, 57774, 57775, 57776, 57777, 57778, 57779, 57780, 
    57781, 57782, 57783, 57784, 57785, 57786, 57787, 57788, 57789, 57790, 
    57791, 57792, 57793, 57794, 57795, 57796, 57797, 57798, 57799, 57800, 
    57801, 57802, 57803, 57804, 57805, 57806, 57807, 57808, 57809, 57810, 
    57811, 57812, 57813, 57814, 57815, 57816, 57817, 57818, 57819, 57820, 
    57821, 57822, 57823, 57824, 57825, 57826, 57827, 57828, 57829, 57830, 
    57831, 57832, 57833, 57834, 57835, 57836, 57837, 57838, 57839, 57840, 
    57841, 57842, 57843, 57844, 57845, 57846, 57847, 57848, 57849, 57850, 
    57851, 57852, 57853, 57854, 57855, 57856, 57857, 57858, 57859, 57860, 
    57861, 57862, 57863, 57864, 57865, 57866, 57867, 57868, 57869, 57870, 
    57871, 57872, 57873, 57874, 57875, 57876, 57877, 57878, 57879, 57880, 
    57881, 57882, 57883, 57884, 57885, 57886, 57887, 57888, 57889, 57890, 
    57891, 57892, 57893, 57894, 57895, 57896, 57897, 57898, 57899, 57900, 
    57901, 57902, 57903, 57904, 57905, 57906, 57907, 57908, 57909, 57910, 
    57911, 57912, 57913, 57914, 57915, 57916, 57917, 57918, 57919, 57920, 
    57921, 57922, 57923, 57924, 57925, 57926, 57927, 57928, 57929, 57930, 
    57931, 57932, 57933, 57934, 57935, 57936, 57937, 57938, 57939, 57940, 
    57941, 57942, 57943, 57944, 57945, 57946, 57947, 57948, 57949, 57950, 
    57951, 57952, 57953, 57954, 57955, 57956, 57957, 57958, 57959, 57960, 
    57961, 57962, 57963, 57964, 57965, 57966, 57967, 57968, 57969, 57970, 
    57971, 57972, 57973, 57974, 57975, 57976, 57977, 57978, 57979, 57980, 
    57981, 57982, 57983, 57984, 57985, 57986, 57987, 57988, 57989, 57990, 
    57991, 57992, 57993, 57994, 57995, 57996, 57997, 57998, 57999, 58000, 
    58001, 58002, 58003, 58004, 58005, 58006, 58007, 58008, 58009, 58010, 
    58011, 58012, 58013, 58014, 58015, 58016, 58017, 58018, 58019, 58020, 
    58021, 58022, 58023, 58024, 58025, 58026, 58027, 58028, 58029, 58030, 
    58031, 58032, 58033, 58034, 58035, 58036, 58037, 58038, 58039, 58040, 
    58041, 58042, 58043, 58044, 58045, 58046, 58047, 58048, 58049, 58050, 
    58051, 58052, 58053, 58054, 58055, 58056, 58057, 58058, 58059, 58060, 
    58061, 58062, 58063, 58064, 58065, 58066, 58067, 58068, 58069, 58070, 
    58071, 58072, 58073, 58074, 58075, 58076, 58077, 58078, 58079, 58080, 
    58081, 58082, 58083, 58084, 58085, 58086, 58087, 58088, 58089, 58090, 
    58091, 58092, 58093, 58094, 58095, 58096, 58097, 58098, 58099, 58100, 
    58101, 58102, 58103, 58104, 58105, 58106, 58107, 58108, 58109, 58110, 
    58111, 58112, 58113, 58114, 58115, 58116, 58117, 58118, 58119, 58120, 
    58121, 58122, 58123, 58124, 58125, 58126, 58127, 58128, 58129, 58130, 
    58131, 58132, 58133, 58134, 58135, 58136, 58137, 58138, 58139, 58140, 
    58141, 58142, 58143, 58144, 58145, 58146, 58147, 58148, 58149, 58150, 
    58151, 58152, 58153, 58154, 58155, 58156, 58157, 58158, 58159, 58160, 
    58161, 58162, 58163, 58164, 58165, 58166, 58167, 58168, 58169, 58170, 
    58171, 58172, 58173, 58174, 58175, 58176, 58177, 58178, 58179, 58180, 
    58181, 58182, 58183, 58184, 58185, 58186, 58187, 58188, 58189, 58190, 
    58191, 58192, 58193, 58194, 58195, 58196, 58197, 58198, 58199, 58200, 
    58201, 58202, 58203, 58204, 58205, 58206, 58207, 58208, 58209, 58210, 
    58211, 58212, 58213, 58214, 58215, 58216, 58217, 58218, 58219, 58220, 
    58221, 58222, 58223, 58224, 58225, 58226, 58227, 58228, 58229, 58230, 
    58231, 58232, 58233, 58234, 58235, 58236, 58237, 58238, 58239, 58240, 
    58241, 58242, 58243, 58244, 58245, 58246, 58247, 58248, 58249, 58250, 
    58251, 58252, 58253, 58254, 58255, 58256, 58257, 58258, 58259, 58260, 
    58261, 58262, 58263, 58264, 58265, 58266, 58267, 58268, 58269, 58270, 
    58271, 58272, 58273, 58274, 58275, 58276, 58277, 58278, 58279, 58280, 
    58281, 58282, 58283, 58284, 58285, 58286, 58287, 58288, 58289, 58290, 
    58291, 58292, 58293, 58294, 58295, 58296, 58297, 58298, 58299, 58300, 
    58301, 58302, 58303, 58304, 58305, 58306, 58307, 58308, 58309, 58310, 
    58311, 58312, 58313, 58314, 58315, 58316, 58317, 58318, 58319, 58320, 
    58321, 58322, 58323, 58324, 58325, 58326, 58327, 58328, 58329, 58330, 
    58331, 58332, 58333, 58334, 58335, 58336, 58337, 58338, 58339, 58340, 
    58341, 58342, 58343, 58344, 58345, 58346, 58347, 58348, 58349, 58350, 
    58351, 58352, 58353, 58354, 58355, 58356, 58357, 58358, 58359, 58360, 
    58361, 58362, 58363, 58364, 58365, 58366, 58367, 58368, 58369, 58370, 
    58371, 58372, 58373, 58374, 58375, 58376, 58377, 58378, 58379, 58380, 
    58381, 58382, 58383, 58384, 58385, 58386, 58387, 58388, 58389, 58390, 
    58391, 58392, 58393, 58394, 58395, 58396, 58397, 58398, 58399, 58400, 
    58401, 58402, 58403, 58404, 58405, 58406, 58407, 58408, 58409, 58410, 
    58411, 58412, 58413, 58414, 58415, 58416, 58417, 58418, 58419, 58420, 
    58421, 58422, 58423, 58424, 58425, 58426, 58427, 58428, 58429, 58430, 
    58431, 58432, 58433, 58434, 58435, 58436, 58437, 58438, 58439, 58440, 
    58441, 58442, 58443, 58444, 58445, 58446, 58447, 58448, 58449, 58450, 
    58451, 58452, 58453, 58454, 58455, 58456, 58457, 58458, 58459, 58460, 
    58461, 58462, 58463, 58464, 58465, 58466, 58467, 58468, 58469, 58470, 
    58471, 58472, 58473, 58474, 58475, 58476, 58477, 58478, 58479, 58480, 
    58481, 58482, 58483, 58484, 58485, 58486, 58487, 58488, 58489, 58490, 
    58491, 58492, 58493, 58494, 58495, 58496, 58497, 58498, 58499, 58500, 
    58501, 58502, 58503, 58504, 58505, 58506, 58507, 58508, 58509, 58510, 
    58511, 58512, 58513, 58514, 58515, 58516, 58517, 58518, 58519, 58520, 
    58521, 58522, 58523, 58524, 58525, 58526, 58527, 58528, 58529, 58530, 
    58531, 58532, 58533, 58534, 58535, 58536, 58537, 58538, 58539, 58540, 
    58541, 58542, 58543, 58544, 58545, 58546, 58547, 58548, 58549, 58550, 
    58551, 58552, 58553, 58554, 58555, 58556, 58557, 58558, 58559, 58560, 
    58561, 58562, 58563, 58564, 58565, 58566, 58567, 58568, 58569, 58570, 
    58571, 58572, 58573, 58574, 58575, 58576, 58577, 58578, 58579, 58580, 
    58581, 58582, 58583, 58584, 58585, 58586, 58587, 58588, 58589, 58590, 
    58591, 58592, 58593, 58594, 58595, 58596, 58597, 58598, 58599, 58600, 
    58601, 58602, 58603, 58604, 58605, 58606, 58607, 58608, 58609, 58610, 
    58611, 58612, 58613, 58614, 58615, 58616, 58617, 58618, 58619, 58620, 
    58621, 58622, 58623, 58624, 58625, 58626, 58627, 58628, 58629, 58630, 
    58631, 58632, 58633, 58634, 58635, 58636, 58637, 58638, 58639, 58640, 
    58641, 58642, 58643, 58644, 58645, 58646, 58647, 58648, 58649, 58650, 
    58651, 58652, 58653, 58654, 58655, 58656, 58657, 58658, 58659, 58660, 
    58661, 58662, 58663, 58664, 58665, 58666, 58667, 58668, 58669, 58670, 
    58671, 58672, 58673, 58674, 58675, 58676, 58677, 58678, 58679, 58680, 
    58681, 58682, 58683, 58684, 58685, 58686, 58687, 58688, 58689, 58690, 
    58691, 58692, 58693, 58694, 58695, 58696, 58697, 58698, 58699, 58700, 
    58701, 58702, 58703, 58704, 58705, 58706, 58707, 58708, 58709, 58710, 
    58711, 58712, 58713, 58714, 58715, 58716, 58717, 58718, 58719, 58720, 
    58721, 58722, 58723, 58724, 58725, 58726, 58727, 58728, 58729, 58730, 
    58731, 58732, 58733, 58734, 58735, 58736, 58737, 58738, 58739, 58740, 
    58741, 58742, 58743, 58744, 58745, 58746, 58747, 58748, 58749, 58750, 
    58751, 58752, 58753, 58754, 58755, 58756, 58757, 58758, 58759, 58760, 
    58761, 58762, 58763, 58764, 58765, 58766, 58767, 58768, 58769, 58770, 
    58771, 58772, 58773, 58774, 58775, 58776, 58777, 58778, 58779, 58780, 
    58781, 58782, 58783, 58784, 58785, 58786, 58787, 58788, 58789, 58790, 
    58791, 58792, 58793, 58794, 58795, 58796, 58797, 58798, 58799, 58800, 
    58801, 58802, 58803, 58804, 58805, 58806, 58807, 58808, 58809, 58810, 
    58811, 58812, 58813, 58814, 58815, 58816, 58817, 58818, 58819, 58820, 
    58821, 58822, 58823, 58824, 58825, 58826, 58827, 58828, 58829, 58830, 
    58831, 58832, 58833, 58834, 58835, 58836, 58837, 58838, 58839, 58840, 
    58841, 58842, 58843, 58844, 58845, 58846, 58847, 58848, 58849, 58850, 
    58851, 58852, 58853, 58854, 58855, 58856, 58857, 58858, 58859, 58860, 
    58861, 58862, 58863, 58864, 58865, 58866, 58867, 58868, 58869, 58870, 
    58871, 58872, 58873, 58874, 58875, 58876, 58877, 58878, 58879, 58880, 
    58881, 58882, 58883, 58884, 58885, 58886, 58887, 58888, 58889, 58890, 
    58891, 58892, 58893, 58894, 58895, 58896, 58897, 58898, 58899, 58900, 
    58901, 58902, 58903, 58904, 58905, 58906, 58907, 58908, 58909, 58910, 
    58911, 58912, 58913, 58914, 58915, 58916, 58917, 58918, 58919, 58920, 
    58921, 58922, 58923, 58924, 58925, 58926, 58927, 58928, 58929, 58930, 
    58931, 58932, 58933, 58934, 58935, 58936, 58937, 58938, 58939, 58940, 
    58941, 58942, 58943, 58944, 58945, 58946, 58947, 58948, 58949, 58950, 
    58951, 58952, 58953, 58954, 58955, 58956, 58957, 58958, 58959, 58960, 
    58961, 58962, 58963, 58964, 58965, 58966, 58967, 58968, 58969, 58970, 
    58971, 58972, 58973, 58974, 58975, 58976, 58977, 58978, 58979, 58980, 
    58981, 58982, 58983, 58984, 58985, 58986, 58987, 58988, 58989, 58990, 
    58991, 58992, 58993, 58994, 58995, 58996, 58997, 58998, 58999, 59000, 
    59001, 59002, 59003, 59004, 59005, 59006, 59007, 59008, 59009, 59010, 
    59011, 59012, 59013, 59014, 59015, 59016, 59017, 59018, 59019, 59020, 
    59021, 59022, 59023, 59024, 59025, 59026, 59027, 59028, 59029, 59030, 
    59031, 59032, 59033, 59034, 59035, 59036, 59037, 59038, 59039, 59040, 
    59041, 59042, 59043, 59044, 59045, 59046, 59047, 59048, 59049, 59050, 
    59051, 59052, 59053, 59054, 59055, 59056, 59057, 59058, 59059, 59060, 
    59061, 59062, 59063, 59064, 59065, 59066, 59067, 59068, 59069, 59070, 
    59071, 59072, 59073, 59074, 59075, 59076, 59077, 59078, 59079, 59080, 
    59081, 59082, 59083, 59084, 59085, 59086, 59087, 59088, 59089, 59090, 
    59091, 59092, 59093, 59094, 59095, 59096, 59097, 59098, 59099, 59100, 
    59101, 59102, 59103, 59104, 59105, 59106, 59107, 59108, 59109, 59110, 
    59111, 59112, 59113, 59114, 59115, 59116, 59117, 59118, 59119, 59120, 
    59121, 59122, 59123, 59124, 59125, 59126, 59127, 59128, 59129, 59130, 
    59131, 59132, 59133, 59134, 59135, 59136, 59137, 59138, 59139, 59140, 
    59141, 59142, 59143, 59144, 59145, 59146, 59147, 59148, 59149, 59150, 
    59151, 59152, 59153, 59154, 59155, 59156, 59157, 59158, 59159, 59160, 
    59161, 59162, 59163, 59164, 59165, 59166, 59167, 59168, 59169, 59170, 
    59171, 59172, 59173, 59174, 59175, 59176, 59177, 59178, 59179, 59180, 
    59181, 59182, 59183, 59184, 59185, 59186, 59187, 59188, 59189, 59190, 
    59191, 59192, 59193, 59194, 59195, 59196, 59197, 59198, 59199, 59200, 
    59201, 59202, 59203, 59204, 59205, 59206, 59207, 59208, 59209, 59210, 
    59211, 59212, 59213, 59214, 59215, 59216, 59217, 59218, 59219, 59220, 
    59221, 59222, 59223, 59224, 59225, 59226, 59227, 59228, 59229, 59230, 
    59231, 59232, 59233, 59234, 59235, 59236, 59237, 59238, 59239, 59240, 
    59241, 59242, 59243, 59244, 59245, 59246, 59247, 59248, 59249, 59250, 
    59251, 59252, 59253, 59254, 59255, 59256, 59257, 59258, 59259, 59260, 
    59261, 59262, 59263, 59264, 59265, 59266, 59267, 59268, 59269, 59270, 
    59271, 59272, 59273, 59274, 59275, 59276, 59277, 59278, 59279, 59280, 
    59281, 59282, 59283, 59284, 59285, 59286, 59287, 59288, 59289, 59290, 
    59291, 59292, 59293, 59294, 59295, 59296, 59297, 59298, 59299, 59300, 
    59301, 59302, 59303, 59304, 59305, 59306, 59307, 59308, 59309, 59310, 
    59311, 59312, 59313, 59314, 59315, 59316, 59317, 59318, 59319, 59320, 
    59321, 59322, 59323, 59324, 59325, 59326, 59327, 59328, 59329, 59330, 
    59331, 59332, 59333, 59334, 59335, 59336, 59337, 59338, 59339, 59340, 
    59341, 59342, 59343, 59344, 59345, 59346, 59347, 59348, 59349, 59350, 
    59351, 59352, 59353, 59354, 59355, 59356, 59357, 59358, 59359, 59360, 
    59361, 59362, 59363, 59364, 59365, 59366, 59367, 59368, 59369, 59370, 
    59371, 59372, 59373, 59374, 59375, 59376, 59377, 59378, 59379, 59380, 
    59381, 59382, 59383, 59384, 59385, 59386, 59387, 59388, 59389, 59390, 
    59391, 59392, 59393, 59394, 59395, 59396, 59397, 59398, 59399, 59400, 
    59401, 59402, 59403, 59404, 59405, 59406, 59407, 59408, 59409, 59410, 
    59411, 59412, 59413, 59414, 59415, 59416, 59417, 59418, 59419, 59420, 
    59421, 59422, 59423, 59424, 59425, 59426, 59427, 59428, 59429, 59430, 
    59431, 59432, 59433, 59434, 59435, 59436, 59437, 59438, 59439, 59440, 
    59441, 59442, 59443, 59444, 59445, 59446, 59447, 59448, 59449, 59450, 
    59451, 59452, 59453, 59454, 59455, 59456, 59457, 59458, 59459, 59460, 
    59461, 59462, 59463, 59464, 59465, 59466, 59467, 59468, 59469, 59470, 
    59471, 59472, 59473, 59474, 59475, 59476, 59477, 59478, 59479, 59480, 
    59481, 59482, 59483, 59484, 59485, 59486, 59487, 59488, 59489, 59490, 
    59491, 59492, 59493, 59494, 59495, 59496, 59497, 59498, 59499, 59500, 
    59501, 59502, 59503, 59504, 59505, 59506, 59507, 59508, 59509, 59510, 
    59511, 59512, 59513, 59514, 59515, 59516, 59517, 59518, 59519, 59520, 
    59521, 59522, 59523, 59524, 59525, 59526, 59527, 59528, 59529, 59530, 
    59531, 59532, 59533, 59534, 59535, 59536, 59537, 59538, 59539, 59540, 
    59541, 59542, 59543, 59544, 59545, 59546, 59547, 59548, 59549, 59550, 
    59551, 59552, 59553, 59554, 59555, 59556, 59557, 59558, 59559, 59560, 
    59561, 59562, 59563, 59564, 59565, 59566, 59567, 59568, 59569, 59570, 
    59571, 59572, 59573, 59574, 59575, 59576, 59577, 59578, 59579, 59580, 
    59581, 59582, 59583, 59584, 59585, 59586, 59587, 59588, 59589, 59590, 
    59591, 59592, 59593, 59594, 59595, 59596, 59597, 59598, 59599, 59600, 
    59601, 59602, 59603, 59604, 59605, 59606, 59607, 59608, 59609, 59610, 
    59611, 59612, 59613, 59614, 59615, 59616, 59617, 59618, 59619, 59620, 
    59621, 59622, 59623, 59624, 59625, 59626, 59627, 59628, 59629, 59630, 
    59631, 59632, 59633, 59634, 59635, 59636, 59637, 59638, 59639, 59640, 
    59641, 59642, 59643, 59644, 59645, 59646, 59647, 59648, 59649, 59650, 
    59651, 59652, 59653, 59654, 59655, 59656, 59657, 59658, 59659, 59660, 
    59661, 59662, 59663, 59664, 59665, 59666, 59667, 59668, 59669, 59670, 
    59671, 59672, 59673, 59674, 59675, 59676, 59677, 59678, 59679, 59680, 
    59681, 59682, 59683, 59684, 59685, 59686, 59687, 59688, 59689, 59690, 
    59691, 59692, 59693, 59694, 59695, 59696, 59697, 59698, 59699, 59700, 
    59701, 59702, 59703, 59704, 59705, 59706, 59707, 59708, 59709, 59710, 
    59711, 59712, 59713, 59714, 59715, 59716, 59717, 59718, 59719, 59720, 
    59721, 59722, 59723, 59724, 59725, 59726, 59727, 59728, 59729, 59730, 
    59731, 59732, 59733, 59734, 59735, 59736, 59737, 59738, 59739, 59740, 
    59741, 59742, 59743, 59744, 59745, 59746, 59747, 59748, 59749, 59750, 
    59751, 59752, 59753, 59754, 59755, 59756, 59757, 59758, 59759, 59760, 
    59761, 59762, 59763, 59764, 59765, 59766, 59767, 59768, 59769, 59770, 
    59771, 59772, 59773, 59774, 59775, 59776, 59777, 59778, 59779, 59780, 
    59781, 59782, 59783, 59784, 59785, 59786, 59787, 59788, 59789, 59790, 
    59791, 59792, 59793, 59794, 59795, 59796, 59797, 59798, 59799, 59800, 
    59801, 59802, 59803, 59804, 59805, 59806, 59807, 59808, 59809, 59810, 
    59811, 59812, 59813, 59814, 59815, 59816, 59817, 59818, 59819, 59820, 
    59821, 59822, 59823, 59824, 59825, 59826, 59827, 59828, 59829, 59830, 
    59831, 59832, 59833, 59834, 59835, 59836, 59837, 59838, 59839, 59840, 
    59841, 59842, 59843, 59844, 59845, 59846, 59847, 59848, 59849, 59850, 
    59851, 59852, 59853, 59854, 59855, 59856, 59857, 59858, 59859, 59860, 
    59861, 59862, 59863, 59864, 59865, 59866, 59867, 59868, 59869, 59870, 
    59871, 59872, 59873, 59874, 59875, 59876, 59877, 59878, 59879, 59880, 
    59881, 59882, 59883, 59884, 59885, 59886, 59887, 59888, 59889, 59890, 
    59891, 59892, 59893, 59894, 59895, 59896, 59897, 59898, 59899, 59900, 
    59901, 59902, 59903, 59904, 59905, 59906, 59907, 59908, 59909, 59910, 
    59911, 59912, 59913, 59914, 59915, 59916, 59917, 59918, 59919, 59920, 
    59921, 59922, 59923, 59924, 59925, 59926, 59927, 59928, 59929, 59930, 
    59931, 59932, 59933, 59934, 59935, 59936, 59937, 59938, 59939, 59940, 
    59941, 59942, 59943, 59944, 59945, 59946, 59947, 59948, 59949, 59950, 
    59951, 59952, 59953, 59954, 59955, 59956, 59957, 59958, 59959, 59960, 
    59961, 59962, 59963, 59964, 59965, 59966, 59967, 59968, 59969, 59970, 
    59971, 59972, 59973, 59974, 59975, 59976, 59977, 59978, 59979, 59980, 
    59981, 59982, 59983, 59984, 59985, 59986, 59987, 59988, 59989, 59990, 
    59991, 59992, 59993, 59994, 59995, 59996, 59997, 59998, 59999, 60000, 
    60001, 60002, 60003, 60004, 60005, 60006, 60007, 60008, 60009, 60010, 
    60011, 60012, 60013, 60014, 60015, 60016, 60017, 60018, 60019, 60020, 
    60021, 60022, 60023, 60024, 60025, 60026, 60027, 60028, 60029, 60030, 
    60031, 60032, 60033, 60034, 60035, 60036, 60037, 60038, 60039, 60040, 
    60041, 60042, 60043, 60044, 60045, 60046, 60047, 60048, 60049, 60050, 
    60051, 60052, 60053, 60054, 60055, 60056, 60057, 60058, 60059, 60060, 
    60061, 60062, 60063, 60064, 60065, 60066, 60067, 60068, 60069, 60070, 
    60071, 60072, 60073, 60074, 60075, 60076, 60077, 60078, 60079, 60080, 
    60081, 60082, 60083, 60084, 60085, 60086, 60087, 60088, 60089, 60090, 
    60091, 60092, 60093, 60094, 60095, 60096, 60097, 60098, 60099, 60100, 
    60101, 60102, 60103, 60104, 60105, 60106, 60107, 60108, 60109, 60110, 
    60111, 60112, 60113, 60114, 60115, 60116, 60117, 60118, 60119, 60120, 
    60121, 60122, 60123, 60124, 60125, 60126, 60127, 60128, 60129, 60130, 
    60131, 60132, 60133, 60134, 60135, 60136, 60137, 60138, 60139, 60140, 
    60141, 60142, 60143, 60144, 60145, 60146, 60147, 60148, 60149, 60150, 
    60151, 60152, 60153, 60154, 60155, 60156, 60157, 60158, 60159, 60160, 
    60161, 60162, 60163, 60164, 60165, 60166, 60167, 60168, 60169, 60170, 
    60171, 60172, 60173, 60174, 60175, 60176, 60177, 60178, 60179, 60180, 
    60181, 60182, 60183, 60184, 60185, 60186, 60187, 60188, 60189, 60190, 
    60191, 60192, 60193, 60194, 60195, 60196, 60197, 60198, 60199, 60200, 
    60201, 60202, 60203, 60204, 60205, 60206, 60207, 60208, 60209, 60210, 
    60211, 60212, 60213, 60214, 60215, 60216, 60217, 60218, 60219, 60220, 
    60221, 60222, 60223, 60224, 60225, 60226, 60227, 60228, 60229, 60230, 
    60231, 60232, 60233, 60234, 60235, 60236, 60237, 60238, 60239, 60240, 
    60241, 60242, 60243, 60244, 60245, 60246, 60247, 60248, 60249, 60250, 
    60251, 60252, 60253, 60254, 60255, 60256, 60257, 60258, 60259, 60260, 
    60261, 60262, 60263, 60264, 60265, 60266, 60267, 60268, 60269, 60270, 
    60271, 60272, 60273, 60274, 60275, 60276, 60277, 60278, 60279, 60280, 
    60281, 60282, 60283, 60284, 60285, 60286, 60287, 60288, 60289, 60290, 
    60291, 60292, 60293, 60294, 60295, 60296, 60297, 60298, 60299, 60300, 
    60301, 60302, 60303, 60304, 60305, 60306, 60307, 60308, 60309, 60310, 
    60311, 60312, 60313, 60314, 60315, 60316, 60317, 60318, 60319, 60320, 
    60321, 60322, 60323, 60324, 60325, 60326, 60327, 60328, 60329, 60330, 
    60331, 60332, 60333, 60334, 60335, 60336, 60337, 60338, 60339, 60340, 
    60341, 60342, 60343, 60344, 60345, 60346, 60347, 60348, 60349, 60350, 
    60351, 60352, 60353, 60354, 60355, 60356, 60357, 60358, 60359, 60360, 
    60361, 60362, 60363, 60364, 60365, 60366, 60367, 60368, 60369, 60370, 
    60371, 60372, 60373, 60374, 60375, 60376, 60377, 60378, 60379, 60380, 
    60381, 60382, 60383, 60384, 60385, 60386, 60387, 60388, 60389, 60390, 
    60391, 60392, 60393, 60394, 60395, 60396, 60397, 60398, 60399, 60400, 
    60401, 60402, 60403, 60404, 60405, 60406, 60407, 60408, 60409, 60410, 
    60411, 60412, 60413, 60414, 60415, 60416, 60417, 60418, 60419, 60420, 
    60421, 60422, 60423, 60424, 60425, 60426, 60427, 60428, 60429, 60430, 
    60431, 60432, 60433, 60434, 60435, 60436, 60437, 60438, 60439, 60440, 
    60441, 60442, 60443, 60444, 60445, 60446, 60447, 60448, 60449, 60450, 
    60451, 60452, 60453, 60454, 60455, 60456, 60457, 60458, 60459, 60460, 
    60461, 60462, 60463, 60464, 60465, 60466, 60467, 60468, 60469, 60470, 
    60471, 60472, 60473, 60474, 60475, 60476, 60477, 60478, 60479, 60480, 
    60481, 60482, 60483, 60484, 60485, 60486, 60487, 60488, 60489, 60490, 
    60491, 60492, 60493, 60494, 60495, 60496, 60497, 60498, 60499, 60500, 
    60501, 60502, 60503, 60504, 60505, 60506, 60507, 60508, 60509, 60510, 
    60511, 60512, 60513, 60514, 60515, 60516, 60517, 60518, 60519, 60520, 
    60521, 60522, 60523, 60524, 60525, 60526, 60527, 60528, 60529, 60530, 
    60531, 60532, 60533, 60534, 60535, 60536, 60537, 60538, 60539, 60540, 
    60541, 60542, 60543, 60544, 60545, 60546, 60547, 60548, 60549, 60550, 
    60551, 60552, 60553, 60554, 60555, 60556, 60557, 60558, 60559, 60560, 
    60561, 60562, 60563, 60564, 60565, 60566, 60567, 60568, 60569, 60570, 
    60571, 60572, 60573, 60574, 60575, 60576, 60577, 60578, 60579, 60580, 
    60581, 60582, 60583, 60584, 60585, 60586, 60587, 60588, 60589, 60590, 
    60591, 60592, 60593, 60594, 60595, 60596, 60597, 60598, 60599, 60600, 
    60601, 60602, 60603, 60604, 60605, 60606, 60607, 60608, 60609, 60610, 
    60611, 60612, 60613, 60614, 60615, 60616, 60617, 60618, 60619, 60620, 
    60621, 60622, 60623, 60624, 60625, 60626, 60627, 60628, 60629, 60630, 
    60631, 60632, 60633, 60634, 60635, 60636, 60637, 60638, 60639, 60640, 
    60641, 60642, 60643, 60644, 60645, 60646, 60647, 60648, 60649, 60650, 
    60651, 60652, 60653, 60654, 60655, 60656, 60657, 60658, 60659, 60660, 
    60661, 60662, 60663, 60664, 60665, 60666, 60667, 60668, 60669, 60670, 
    60671, 60672, 60673, 60674, 60675, 60676, 60677, 60678, 60679, 60680, 
    60681, 60682, 60683, 60684, 60685, 60686, 60687, 60688, 60689, 60690, 
    60691, 60692, 60693, 60694, 60695, 60696, 60697, 60698, 60699, 60700, 
    60701, 60702, 60703, 60704, 60705, 60706, 60707, 60708, 60709, 60710, 
    60711, 60712, 60713, 60714, 60715, 60716, 60717, 60718, 60719, 60720, 
    60721, 60722, 60723, 60724, 60725, 60726, 60727, 60728, 60729, 60730, 
    60731, 60732, 60733, 60734, 60735, 60736, 60737, 60738, 60739, 60740, 
    60741, 60742, 60743, 60744, 60745, 60746, 60747, 60748, 60749, 60750, 
    60751, 60752, 60753, 60754, 60755, 60756, 60757, 60758, 60759, 60760, 
    60761, 60762, 60763, 60764, 60765, 60766, 60767, 60768, 60769, 60770, 
    60771, 60772, 60773, 60774, 60775, 60776, 60777, 60778, 60779, 60780, 
    60781, 60782, 60783, 60784, 60785, 60786, 60787, 60788, 60789, 60790, 
    60791, 60792, 60793, 60794, 60795, 60796, 60797, 60798, 60799, 60800, 
    60801, 60802, 60803, 60804, 60805, 60806, 60807, 60808, 60809, 60810, 
    60811, 60812, 60813, 60814, 60815, 60816, 60817, 60818, 60819, 60820, 
    60821, 60822, 60823, 60824, 60825, 60826, 60827, 60828, 60829, 60830, 
    60831, 60832, 60833, 60834, 60835, 60836, 60837, 60838, 60839, 60840, 
    60841, 60842, 60843, 60844, 60845, 60846, 60847, 60848, 60849, 60850, 
    60851, 60852, 60853, 60854, 60855, 60856, 60857, 60858, 60859, 60860, 
    60861, 60862, 60863, 60864, 60865, 60866, 60867, 60868, 60869, 60870, 
    60871, 60872, 60873, 60874, 60875, 60876, 60877, 60878, 60879, 60880, 
    60881, 60882, 60883, 60884, 60885, 60886, 60887, 60888, 60889, 60890, 
    60891, 60892, 60893, 60894, 60895, 60896, 60897, 60898, 60899, 60900, 
    60901, 60902, 60903, 60904, 60905, 60906, 60907, 60908, 60909, 60910, 
    60911, 60912, 60913, 60914, 60915, 60916, 60917, 60918, 60919, 60920, 
    60921, 60922, 60923, 60924, 60925, 60926, 60927, 60928, 60929, 60930, 
    60931, 60932, 60933, 60934, 60935, 60936, 60937, 60938, 60939, 60940, 
    60941, 60942, 60943, 60944, 60945, 60946, 60947, 60948, 60949, 60950, 
    60951, 60952, 60953, 60954, 60955, 60956, 60957, 60958, 60959, 60960, 
    60961, 60962, 60963, 60964, 60965, 60966, 60967, 60968, 60969, 60970, 
    60971, 60972, 60973, 60974, 60975, 60976, 60977, 60978, 60979, 60980, 
    60981, 60982, 60983, 60984, 60985, 60986, 60987, 60988, 60989, 60990, 
    60991, 60992, 60993, 60994, 60995, 60996, 60997, 60998, 60999, 61000, 
    61001, 61002, 61003, 61004, 61005, 61006, 61007, 61008, 61009, 61010, 
    61011, 61012, 61013, 61014, 61015, 61016, 61017, 61018, 61019, 61020, 
    61021, 61022, 61023, 61024, 61025, 61026, 61027, 61028, 61029, 61030, 
    61031, 61032, 61033, 61034, 61035, 61036, 61037, 61038, 61039, 61040, 
    61041, 61042, 61043, 61044, 61045, 61046, 61047, 61048, 61049, 61050, 
    61051, 61052, 61053, 61054, 61055, 61056, 61057, 61058, 61059, 61060, 
    61061, 61062, 61063, 61064, 61065, 61066, 61067, 61068, 61069, 61070, 
    61071, 61072, 61073, 61074, 61075, 61076, 61077, 61078, 61079, 61080, 
    61081, 61082, 61083, 61084, 61085, 61086, 61087, 61088, 61089, 61090, 
    61091, 61092, 61093, 61094, 61095, 61096, 61097, 61098, 61099, 61100, 
    61101, 61102, 61103, 61104, 61105, 61106, 61107, 61108, 61109, 61110, 
    61111, 61112, 61113, 61114, 61115, 61116, 61117, 61118, 61119, 61120, 
    61121, 61122, 61123, 61124, 61125, 61126, 61127, 61128, 61129, 61130, 
    61131, 61132, 61133, 61134, 61135, 61136, 61137, 61138, 61139, 61140, 
    61141, 61142, 61143, 61144, 61145, 61146, 61147, 61148, 61149, 61150, 
    61151, 61152, 61153, 61154, 61155, 61156, 61157, 61158, 61159, 61160, 
    61161, 61162, 61163, 61164, 61165, 61166, 61167, 61168, 61169, 61170, 
    61171, 61172, 61173, 61174, 61175, 61176, 61177, 61178, 61179, 61180, 
    61181, 61182, 61183, 61184, 61185, 61186, 61187, 61188, 61189, 61190, 
    61191, 61192, 61193, 61194, 61195, 61196, 61197, 61198, 61199, 61200, 
    61201, 61202, 61203, 61204, 61205, 61206, 61207, 61208, 61209, 61210, 
    61211, 61212, 61213, 61214, 61215, 61216, 61217, 61218, 61219, 61220, 
    61221, 61222, 61223, 61224, 61225, 61226, 61227, 61228, 61229, 61230, 
    61231, 61232, 61233, 61234, 61235, 61236, 61237, 61238, 61239, 61240, 
    61241, 61242, 61243, 61244, 61245, 61246, 61247, 61248, 61249, 61250, 
    61251, 61252, 61253, 61254, 61255, 61256, 61257, 61258, 61259, 61260, 
    61261, 61262, 61263, 61264, 61265, 61266, 61267, 61268, 61269, 61270, 
    61271, 61272, 61273, 61274, 61275, 61276, 61277, 61278, 61279, 61280, 
    61281, 61282, 61283, 61284, 61285, 61286, 61287, 61288, 61289, 61290, 
    61291, 61292, 61293, 61294, 61295, 61296, 61297, 61298, 61299, 61300, 
    61301, 61302, 61303, 61304, 61305, 61306, 61307, 61308, 61309, 61310, 
    61311, 61312, 61313, 61314, 61315, 61316, 61317, 61318, 61319, 61320, 
    61321, 61322, 61323, 61324, 61325, 61326, 61327, 61328, 61329, 61330, 
    61331, 61332, 61333, 61334, 61335, 61336, 61337, 61338, 61339, 61340, 
    61341, 61342, 61343, 61344, 61345, 61346, 61347, 61348, 61349, 61350, 
    61351, 61352, 61353, 61354, 61355, 61356, 61357, 61358, 61359, 61360, 
    61361, 61362, 61363, 61364, 61365, 61366, 61367, 61368, 61369, 61370, 
    61371, 61372, 61373, 61374, 61375, 61376, 61377, 61378, 61379, 61380, 
    61381, 61382, 61383, 61384, 61385, 61386, 61387, 61388, 61389, 61390, 
    61391, 61392, 61393, 61394, 61395, 61396, 61397, 61398, 61399, 61400, 
    61401, 61402, 61403, 61404, 61405, 61406, 61407, 61408, 61409, 61410, 
    61411, 61412, 61413, 61414, 61415, 61416, 61417, 61418, 61419, 61420, 
    61421, 61422, 61423, 61424, 61425, 61426, 61427, 61428, 61429, 61430, 
    61431, 61432, 61433, 61434, 61435, 61436, 61437, 61438, 61439, 61440, 
    61441, 61442, 61443, 61444, 61445, 61446, 61447, 61448, 61449, 61450, 
    61451, 61452, 61453, 61454, 61455, 61456, 61457, 61458, 61459, 61460, 
    61461, 61462, 61463, 61464, 61465, 61466, 61467, 61468, 61469, 61470, 
    61471, 61472, 61473, 61474, 61475, 61476, 61477, 61478, 61479, 61480, 
    61481, 61482, 61483, 61484, 61485, 61486, 61487, 61488, 61489, 61490, 
    61491, 61492, 61493, 61494, 61495, 61496, 61497, 61498, 61499, 61500, 
    61501, 61502, 61503, 61504, 61505, 61506, 61507, 61508, 61509, 61510, 
    61511, 61512, 61513, 61514, 61515, 61516, 61517, 61518, 61519, 61520, 
    61521, 61522, 61523, 61524, 61525, 61526, 61527, 61528, 61529, 61530, 
    61531, 61532, 61533, 61534, 61535, 61536, 61537, 61538, 61539, 61540, 
    61541, 61542, 61543, 61544, 61545, 61546, 61547, 61548, 61549, 61550, 
    61551, 61552, 61553, 61554, 61555, 61556, 61557, 61558, 61559, 61560, 
    61561, 61562, 61563, 61564, 61565, 61566, 61567, 61568, 61569, 61570, 
    61571, 61572, 61573, 61574, 61575, 61576, 61577, 61578, 61579, 61580, 
    61581, 61582, 61583, 61584, 61585, 61586, 61587, 61588, 61589, 61590, 
    61591, 61592, 61593, 61594, 61595, 61596, 61597, 61598, 61599, 61600, 
    61601, 61602, 61603, 61604, 61605, 61606, 61607, 61608, 61609, 61610, 
    61611, 61612, 61613, 61614, 61615, 61616, 61617, 61618, 61619, 61620, 
    61621, 61622, 61623, 61624, 61625, 61626, 61627, 61628, 61629, 61630, 
    61631, 61632, 61633, 61634, 61635, 61636, 61637, 61638, 61639, 61640, 
    61641, 61642, 61643, 61644, 61645, 61646, 61647, 61648, 61649, 61650, 
    61651, 61652, 61653, 61654, 61655, 61656, 61657, 61658, 61659, 61660, 
    61661, 61662, 61663, 61664, 61665, 61666, 61667, 61668, 61669, 61670, 
    61671, 61672, 61673, 61674, 61675, 61676, 61677, 61678, 61679, 61680, 
    61681, 61682, 61683, 61684, 61685, 61686, 61687, 61688, 61689, 61690, 
    61691, 61692, 61693, 61694, 61695, 61696, 61697, 61698, 61699, 61700, 
    61701, 61702, 61703, 61704, 61705, 61706, 61707, 61708, 61709, 61710, 
    61711, 61712, 61713, 61714, 61715, 61716, 61717, 61718, 61719, 61720, 
    61721, 61722, 61723, 61724, 61725, 61726, 61727, 61728, 61729, 61730, 
    61731, 61732, 61733, 61734, 61735, 61736, 61737, 61738, 61739, 61740, 
    61741, 61742, 61743, 61744, 61745, 61746, 61747, 61748, 61749, 61750, 
    61751, 61752, 61753, 61754, 61755, 61756, 61757, 61758, 61759, 61760, 
    61761, 61762, 61763, 61764, 61765, 61766, 61767, 61768, 61769, 61770, 
    61771, 61772, 61773, 61774, 61775, 61776, 61777, 61778, 61779, 61780, 
    61781, 61782, 61783, 61784, 61785, 61786, 61787, 61788, 61789, 61790, 
    61791, 61792, 61793, 61794, 61795, 61796, 61797, 61798, 61799, 61800, 
    61801, 61802, 61803, 61804, 61805, 61806, 61807, 61808, 61809, 61810, 
    61811, 61812, 61813, 61814, 61815, 61816, 61817, 61818, 61819, 61820, 
    61821, 61822, 61823, 61824, 61825, 61826, 61827, 61828, 61829, 61830, 
    61831, 61832, 61833, 61834, 61835, 61836, 61837, 61838, 61839, 61840, 
    61841, 61842, 61843, 61844, 61845, 61846, 61847, 61848, 61849, 61850, 
    61851, 61852, 61853, 61854, 61855, 61856, 61857, 61858, 61859, 61860, 
    61861, 61862, 61863, 61864, 61865, 61866, 61867, 61868, 61869, 61870, 
    61871, 61872, 61873, 61874, 61875, 61876, 61877, 61878, 61879, 61880, 
    61881, 61882, 61883, 61884, 61885, 61886, 61887, 61888, 61889, 61890, 
    61891, 61892, 61893, 61894, 61895, 61896, 61897, 61898, 61899, 61900, 
    61901, 61902, 61903, 61904, 61905, 61906, 61907, 61908, 61909, 61910, 
    61911, 61912, 61913, 61914, 61915, 61916, 61917, 61918, 61919, 61920, 
    61921, 61922, 61923, 61924, 61925, 61926, 61927, 61928, 61929, 61930, 
    61931, 61932, 61933, 61934, 61935, 61936, 61937, 61938, 61939, 61940, 
    61941, 61942, 61943, 61944, 61945, 61946, 61947, 61948, 61949, 61950, 
    61951, 61952, 61953, 61954, 61955, 61956, 61957, 61958, 61959, 61960, 
    61961, 61962, 61963, 61964, 61965, 61966, 61967, 61968, 61969, 61970, 
    61971, 61972, 61973, 61974, 61975, 61976, 61977, 61978, 61979, 61980, 
    61981, 61982, 61983, 61984, 61985, 61986, 61987, 61988, 61989, 61990, 
    61991, 61992, 61993, 61994, 61995, 61996, 61997, 61998, 61999, 62000, 
    62001, 62002, 62003, 62004, 62005, 62006, 62007, 62008, 62009, 62010, 
    62011, 62012, 62013, 62014, 62015, 62016, 62017, 62018, 62019, 62020, 
    62021, 62022, 62023, 62024, 62025, 62026, 62027, 62028, 62029, 62030, 
    62031, 62032, 62033, 62034, 62035, 62036, 62037, 62038, 62039, 62040, 
    62041, 62042, 62043, 62044, 62045, 62046, 62047, 62048, 62049, 62050, 
    62051, 62052, 62053, 62054, 62055, 62056, 62057, 62058, 62059, 62060, 
    62061, 62062, 62063, 62064, 62065, 62066, 62067, 62068, 62069, 62070, 
    62071, 62072, 62073, 62074, 62075, 62076, 62077, 62078, 62079, 62080, 
    62081, 62082, 62083, 62084, 62085, 62086, 62087, 62088, 62089, 62090, 
    62091, 62092, 62093, 62094, 62095, 62096, 62097, 62098, 62099, 62100, 
    62101, 62102, 62103, 62104, 62105, 62106, 62107, 62108, 62109, 62110, 
    62111, 62112, 62113, 62114, 62115, 62116, 62117, 62118, 62119, 62120, 
    62121, 62122, 62123, 62124, 62125, 62126, 62127, 62128, 62129, 62130, 
    62131, 62132, 62133, 62134, 62135, 62136, 62137, 62138, 62139, 62140, 
    62141, 62142, 62143, 62144, 62145, 62146, 62147, 62148, 62149, 62150, 
    62151, 62152, 62153, 62154, 62155, 62156, 62157, 62158, 62159, 62160, 
    62161, 62162, 62163, 62164, 62165, 62166, 62167, 62168, 62169, 62170, 
    62171, 62172, 62173, 62174, 62175, 62176, 62177, 62178, 62179, 62180, 
    62181, 62182, 62183, 62184, 62185, 62186, 62187, 62188, 62189, 62190, 
    62191, 62192, 62193, 62194, 62195, 62196, 62197, 62198, 62199, 62200, 
    62201, 62202, 62203, 62204, 62205, 62206, 62207, 62208, 62209, 62210, 
    62211, 62212, 62213, 62214, 62215, 62216, 62217, 62218, 62219, 62220, 
    62221, 62222, 62223, 62224, 62225, 62226, 62227, 62228, 62229, 62230, 
    62231, 62232, 62233, 62234, 62235, 62236, 62237, 62238, 62239, 62240, 
    62241, 62242, 62243, 62244, 62245, 62246, 62247, 62248, 62249, 62250, 
    62251, 62252, 62253, 62254, 62255, 62256, 62257, 62258, 62259, 62260, 
    62261, 62262, 62263, 62264, 62265, 62266, 62267, 62268, 62269, 62270, 
    62271, 62272, 62273, 62274, 62275, 62276, 62277, 62278, 62279, 62280, 
    62281, 62282, 62283, 62284, 62285, 62286, 62287, 62288, 62289, 62290, 
    62291, 62292, 62293, 62294, 62295, 62296, 62297, 62298, 62299, 62300, 
    62301, 62302, 62303, 62304, 62305, 62306, 62307, 62308, 62309, 62310, 
    62311, 62312, 62313, 62314, 62315, 62316, 62317, 62318, 62319, 62320, 
    62321, 62322, 62323, 62324, 62325, 62326, 62327, 62328, 62329, 62330, 
    62331, 62332, 62333, 62334, 62335, 62336, 62337, 62338, 62339, 62340, 
    62341, 62342, 62343, 62344, 62345, 62346, 62347, 62348, 62349, 62350, 
    62351, 62352, 62353, 62354, 62355, 62356, 62357, 62358, 62359, 62360, 
    62361, 62362, 62363, 62364, 62365, 62366, 62367, 62368, 62369, 62370, 
    62371, 62372, 62373, 62374, 62375, 62376, 62377, 62378, 62379, 62380, 
    62381, 62382, 62383, 62384, 62385, 62386, 62387, 62388, 62389, 62390, 
    62391, 62392, 62393, 62394, 62395, 62396, 62397, 62398, 62399, 62400, 
    62401, 62402, 62403, 62404, 62405, 62406, 62407, 62408, 62409, 62410, 
    62411, 62412, 62413, 62414, 62415, 62416, 62417, 62418, 62419, 62420, 
    62421, 62422, 62423, 62424, 62425, 62426, 62427, 62428, 62429, 62430, 
    62431, 62432, 62433, 62434, 62435, 62436, 62437, 62438, 62439, 62440, 
    62441, 62442, 62443, 62444, 62445, 62446, 62447, 62448, 62449, 62450, 
    62451, 62452, 62453, 62454, 62455, 62456, 62457, 62458, 62459, 62460, 
    62461, 62462, 62463, 62464, 62465, 62466, 62467, 62468, 62469, 62470, 
    62471, 62472, 62473, 62474, 62475, 62476, 62477, 62478, 62479, 62480, 
    62481, 62482, 62483, 62484, 62485, 62486, 62487, 62488, 62489, 62490, 
    62491, 62492, 62493, 62494, 62495, 62496, 62497, 62498, 62499, 62500, 
    62501, 62502, 62503, 62504, 62505, 62506, 62507, 62508, 62509, 62510, 
    62511, 62512, 62513, 62514, 62515, 62516, 62517, 62518, 62519, 62520, 
    62521, 62522, 62523, 62524, 62525, 62526, 62527, 62528, 62529, 62530, 
    62531, 62532, 62533, 62534, 62535, 62536, 62537, 62538, 62539, 62540, 
    62541, 62542, 62543, 62544, 62545, 62546, 62547, 62548, 62549, 62550, 
    62551, 62552, 62553, 62554, 62555, 62556, 62557, 62558, 62559, 62560, 
    62561, 62562, 62563, 62564, 62565, 62566, 62567, 62568, 62569, 62570, 
    62571, 62572, 62573, 62574, 62575, 62576, 62577, 62578, 62579, 62580, 
    62581, 62582, 62583, 62584, 62585, 62586, 62587, 62588, 62589, 62590, 
    62591, 62592, 62593, 62594, 62595, 62596, 62597, 62598, 62599, 62600, 
    62601, 62602, 62603, 62604, 62605, 62606, 62607, 62608, 62609, 62610, 
    62611, 62612, 62613, 62614, 62615, 62616, 62617, 62618, 62619, 62620, 
    62621, 62622, 62623, 62624, 62625, 62626, 62627, 62628, 62629, 62630, 
    62631, 62632, 62633, 62634, 62635, 62636, 62637, 62638, 62639, 62640, 
    62641, 62642, 62643, 62644, 62645, 62646, 62647, 62648, 62649, 62650, 
    62651, 62652, 62653, 62654, 62655, 62656, 62657, 62658, 62659, 62660, 
    62661, 62662, 62663, 62664, 62665, 62666, 62667, 62668, 62669, 62670, 
    62671, 62672, 62673, 62674, 62675, 62676, 62677, 62678, 62679, 62680, 
    62681, 62682, 62683, 62684, 62685, 62686, 62687, 62688, 62689, 62690, 
    62691, 62692, 62693, 62694, 62695, 62696, 62697, 62698, 62699, 62700, 
    62701, 62702, 62703, 62704, 62705, 62706, 62707, 62708, 62709, 62710, 
    62711, 62712, 62713, 62714, 62715, 62716, 62717, 62718, 62719, 62720, 
    62721, 62722, 62723, 62724, 62725, 62726, 62727, 62728, 62729, 62730, 
    62731, 62732, 62733, 62734, 62735, 62736, 62737, 62738, 62739, 62740, 
    62741, 62742, 62743, 62744, 62745, 62746, 62747, 62748, 62749, 62750, 
    62751, 62752, 62753, 62754, 62755, 62756, 62757, 62758, 62759, 62760, 
    62761, 62762, 62763, 62764, 62765, 62766, 62767, 62768, 62769, 62770, 
    62771, 62772, 62773, 62774, 62775, 62776, 62777, 62778, 62779, 62780, 
    62781, 62782, 62783, 62784, 62785, 62786, 62787, 62788, 62789, 62790, 
    62791, 62792, 62793, 62794, 62795, 62796, 62797, 62798, 62799, 62800, 
    62801, 62802, 62803, 62804, 62805, 62806, 62807, 62808, 62809, 62810, 
    62811, 62812, 62813, 62814, 62815, 62816, 62817, 62818, 62819, 62820, 
    62821, 62822, 62823, 62824, 62825, 62826, 62827, 62828, 62829, 62830, 
    62831, 62832, 62833, 62834, 62835, 62836, 62837, 62838, 62839, 62840, 
    62841, 62842, 62843, 62844, 62845, 62846, 62847, 62848, 62849, 62850, 
    62851, 62852, 62853, 62854, 62855, 62856, 62857, 62858, 62859, 62860, 
    62861, 62862, 62863, 62864, 62865, 62866, 62867, 62868, 62869, 62870, 
    62871, 62872, 62873, 62874, 62875, 62876, 62877, 62878, 62879, 62880, 
    62881, 62882, 62883, 62884, 62885, 62886, 62887, 62888, 62889, 62890, 
    62891, 62892, 62893, 62894, 62895, 62896, 62897, 62898, 62899, 62900, 
    62901, 62902, 62903, 62904, 62905, 62906, 62907, 62908, 62909, 62910, 
    62911, 62912, 62913, 62914, 62915, 62916, 62917, 62918, 62919, 62920, 
    62921, 62922, 62923, 62924, 62925, 62926, 62927, 62928, 62929, 62930, 
    62931, 62932, 62933, 62934, 62935, 62936, 62937, 62938, 62939, 62940, 
    62941, 62942, 62943, 62944, 62945, 62946, 62947, 62948, 62949, 62950, 
    62951, 62952, 62953, 62954, 62955, 62956, 62957, 62958, 62959, 62960, 
    62961, 62962, 62963, 62964, 62965, 62966, 62967, 62968, 62969, 62970, 
    62971, 62972, 62973, 62974, 62975, 62976, 62977, 62978, 62979, 62980, 
    62981, 62982, 62983, 62984, 62985, 62986, 62987, 62988, 62989, 62990, 
    62991, 62992, 62993, 62994, 62995, 62996, 62997, 62998, 62999, 63000, 
    63001, 63002, 63003, 63004, 63005, 63006, 63007, 63008, 63009, 63010, 
    63011, 63012, 63013, 63014, 63015, 63016, 63017, 63018, 63019, 63020, 
    63021, 63022, 63023, 63024, 63025, 63026, 63027, 63028, 63029, 63030, 
    63031, 63032, 63033, 63034, 63035, 63036, 63037, 63038, 63039, 63040, 
    63041, 63042, 63043, 63044, 63045, 63046, 63047, 63048, 63049, 63050, 
    63051, 63052, 63053, 63054, 63055, 63056, 63057, 63058, 63059, 63060, 
    63061, 63062, 63063, 63064, 63065, 63066, 63067, 63068, 63069, 63070, 
    63071, 63072, 63073, 63074, 63075, 63076, 63077, 63078, 63079, 63080, 
    63081, 63082, 63083, 63084, 63085, 63086, 63087, 63088, 63089, 63090, 
    63091, 63092, 63093, 63094, 63095, 63096, 63097, 63098, 63099, 63100, 
    63101, 63102, 63103, 63104, 63105, 63106, 63107, 63108, 63109, 63110, 
    63111, 63112, 63113, 63114, 63115, 63116, 63117, 63118, 63119, 63120, 
    63121, 63122, 63123, 63124, 63125, 63126, 63127, 63128, 63129, 63130, 
    63131, 63132, 63133, 63134, 63135, 63136, 63137, 63138, 63139, 63140, 
    63141, 63142, 63143, 63144, 63145, 63146, 63147, 63148, 63149, 63150, 
    63151, 63152, 63153, 63154, 63155, 63156, 63157, 63158, 63159, 63160, 
    63161, 63162, 63163, 63164, 63165, 63166, 63167, 63168, 63169, 63170, 
    63171, 63172, 63173, 63174, 63175, 63176, 63177, 63178, 63179, 63180, 
    63181, 63182, 63183, 63184, 63185, 63186, 63187, 63188, 63189, 63190, 
    63191, 63192, 63193, 63194, 63195, 63196, 63197, 63198, 63199, 63200, 
    63201, 63202, 63203, 63204, 63205, 63206, 63207, 63208, 63209, 63210, 
    63211, 63212, 63213, 63214, 63215, 63216, 63217, 63218, 63219, 63220, 
    63221, 63222, 63223, 63224, 63225, 63226, 63227, 63228, 63229, 63230, 
    63231, 63232, 63233, 63234, 63235, 63236, 63237, 63238, 63239, 63240, 
    63241, 63242, 63243, 63244, 63245, 63246, 63247, 63248, 63249, 63250, 
    63251, 63252, 63253, 63254, 63255, 63256, 63257, 63258, 63259, 63260, 
    63261, 63262, 63263, 63264, 63265, 63266, 63267, 63268, 63269, 63270, 
    63271, 63272, 63273, 63274, 63275, 63276, 63277, 63278, 63279, 63280, 
    63281, 63282, 63283, 63284, 63285, 63286, 63287, 63288, 63289, 63290, 
    63291, 63292, 63293, 63294, 63295, 63296, 63297, 63298, 63299, 63300, 
    63301, 63302, 63303, 63304, 63305, 63306, 63307, 63308, 63309, 63310, 
    63311, 63312, 63313, 63314, 63315, 63316, 63317, 63318, 63319, 63320, 
    63321, 63322, 63323, 63324, 63325, 63326, 63327, 63328, 63329, 63330, 
    63331, 63332, 63333, 63334, 63335, 63336, 63337, 63338, 63339, 63340, 
    63341, 63342, 63343, 63344, 63345, 63346, 63347, 63348, 63349, 63350, 
    63351, 63352, 63353, 63354, 63355, 63356, 63357, 63358, 63359, 63360, 
    63361, 63362, 63363, 63364, 63365, 63366, 63367, 63368, 63369, 63370, 
    63371, 63372, 63373, 63374, 63375, 63376, 63377, 63378, 63379, 63380, 
    63381, 63382, 63383, 63384, 63385, 63386, 63387, 63388, 63389, 63390, 
    63391, 63392, 63393, 63394, 63395, 63396, 63397, 63398, 63399, 63400, 
    63401, 63402, 63403, 63404, 63405, 63406, 63407, 63408, 63409, 63410, 
    63411, 63412, 63413, 63414, 63415, 63416, 63417, 63418, 63419, 63420, 
    63421, 63422, 63423, 63424, 63425, 63426, 63427, 63428, 63429, 63430, 
    63431, 63432, 63433, 63434, 63435, 63436, 63437, 63438, 63439, 63440, 
    63441, 63442, 63443, 63444, 63445, 63446, 63447, 63448, 63449, 63450, 
    63451, 63452, 63453, 63454, 63455, 63456, 63457, 63458, 63459, 63460, 
    63461, 63462, 63463, 63464, 63465, 63466, 63467, 63468, 63469, 63470, 
    63471, 63472, 63473, 63474, 63475, 63476, 63477, 63478, 63479, 63480, 
    63481, 63482, 63483, 63484, 63485, 63486, 63487, 63488, 63489, 63490, 
    63491, 63492, 63493, 63494, 63495, 63496, 63497, 63498, 63499, 63500, 
    63501, 63502, 63503, 63504, 63505, 63506, 63507, 63508, 63509, 63510, 
    63511, 63512, 63513, 63514, 63515, 63516, 63517, 63518, 63519, 63520, 
    63521, 63522, 63523, 63524, 63525, 63526, 63527, 63528, 63529, 63530, 
    63531, 63532, 63533, 63534, 63535, 63536, 63537, 63538, 63539, 63540, 
    63541, 63542, 63543, 63544, 63545, 63546, 63547, 63548, 63549, 63550, 
    63551, 63552, 63553, 63554, 63555, 63556, 63557, 63558, 63559, 63560, 
    63561, 63562, 63563, 63564, 63565, 63566, 63567, 63568, 63569, 63570, 
    63571, 63572, 63573, 63574, 63575, 63576, 63577, 63578, 63579, 63580, 
    63581, 63582, 63583, 63584, 63585, 63586, 63587, 63588, 63589, 63590, 
    63591, 63592, 63593, 63594, 63595, 63596, 63597, 63598, 63599, 63600, 
    63601, 63602, 63603, 63604, 63605, 63606, 63607, 63608, 63609, 63610, 
    63611, 63612, 63613, 63614, 63615, 63616, 63617, 63618, 63619, 63620, 
    63621, 63622, 63623, 63624, 63625, 63626, 63627, 63628, 63629, 63630, 
    63631, 63632, 63633, 63634, 63635, 63636, 63637, 63638, 63639, 63640, 
    63641, 63642, 63643, 63644, 63645, 63646, 63647, 63648, 63649, 63650, 
    63651, 63652, 63653, 63654, 63655, 63656, 63657, 63658, 63659, 63660, 
    63661, 63662, 63663, 63664, 63665, 63666, 63667, 63668, 63669, 63670, 
    63671, 63672, 63673, 63674, 63675, 63676, 63677, 63678, 63679, 63680, 
    63681, 63682, 63683, 63684, 63685, 63686, 63687, 63688, 63689, 63690, 
    63691, 63692, 63693, 63694, 63695, 63696, 63697, 63698, 63699, 63700, 
    63701, 63702, 63703, 63704, 63705, 63706, 63707, 63708, 63709, 63710, 
    63711, 63712, 63713, 63714, 63715, 63716, 63717, 63718, 63719, 63720, 
    63721, 63722, 63723, 63724, 63725, 63726, 63727, 63728, 63729, 63730, 
    63731, 63732, 63733, 63734, 63735, 63736, 63737, 63738, 63739, 63740, 
    63741, 63742, 63743, 63744, 63745, 63746, 63747, 63748, 63749, 63750, 
    63751, 63752, 63753, 63754, 63755, 63756, 63757, 63758, 63759, 63760, 
    63761, 63762, 63763, 63764, 63765, 63766, 63767, 63768, 63769, 63770, 
    63771, 63772, 63773, 63774, 63775, 63776, 63777, 63778, 63779, 63780, 
    63781, 63782, 63783, 63784, 63785, 63786, 63787, 63788, 63789, 63790, 
    63791, 63792, 63793, 63794, 63795, 63796, 63797, 63798, 63799, 63800, 
    63801, 63802, 63803, 63804, 63805, 63806, 63807, 63808, 63809, 63810, 
    63811, 63812, 63813, 63814, 63815, 63816, 63817, 63818, 63819, 63820, 
    63821, 63822, 63823, 63824, 63825, 63826, 63827, 63828, 63829, 63830, 
    63831, 63832, 63833, 63834, 63835, 63836, 63837, 63838, 63839, 63840, 
    63841, 63842, 63843, 63844, 63845, 63846, 63847, 63848, 63849, 63850, 
    63851, 63852, 63853, 63854, 63855, 63856, 63857, 63858, 63859, 63860, 
    63861, 63862, 63863, 63864, 63865, 63866, 63867, 63868, 63869, 63870, 
    63871, 63872, 63873, 63874, 63875, 63876, 63877, 63878, 63879, 63880, 
    63881, 63882, 63883, 63884, 63885, 63886, 63887, 63888, 63889, 63890, 
    63891, 63892, 63893, 63894, 63895, 63896, 63897, 63898, 63899, 63900, 
    63901, 63902, 63903, 63904, 63905, 63906, 63907, 63908, 63909, 63910, 
    63911, 63912, 63913, 63914, 63915, 63916, 63917, 63918, 63919, 63920, 
    63921, 63922, 63923, 63924, 63925, 63926, 63927, 63928, 63929, 63930, 
    63931, 63932, 63933, 63934, 63935, 63936, 63937, 63938, 63939, 63940, 
    63941, 63942, 63943, 63944, 63945, 63946, 63947, 63948, 63949, 63950, 
    63951, 63952, 63953, 63954, 63955, 63956, 63957, 63958, 63959, 63960, 
    63961, 63962, 63963, 63964, 63965, 63966, 63967, 63968, 63969, 63970, 
    63971, 63972, 63973, 63974, 63975, 63976, 63977, 63978, 63979, 63980, 
    63981, 63982, 63983, 63984, 63985, 63986, 63987, 63988, 63989, 63990, 
    63991, 63992, 63993, 63994, 63995, 63996, 63997, 63998, 63999, 64000, 
    64001, 64002, 64003, 64004, 64005, 64006, 64007, 64008, 64009, 64010, 
    64011, 64012, 64013, 64014, 64015, 64016, 64017, 64018, 64019, 64020, 
    64021, 64022, 64023, 64024, 64025, 64026, 64027, 64028, 64029, 64030, 
    64031, 64032, 64033, 64034, 64035, 64036, 64037, 64038, 64039, 64040, 
    64041, 64042, 64043, 64044, 64045, 64046, 64047, 64048, 64049, 64050, 
    64051, 64052, 64053, 64054, 64055, 64056, 64057, 64058, 64059, 64060, 
    64061, 64062, 64063, 64064, 64065, 64066, 64067, 64068, 64069, 64070, 
    64071, 64072, 64073, 64074, 64075, 64076, 64077, 64078, 64079, 64080, 
    64081, 64082, 64083, 64084, 64085, 64086, 64087, 64088, 64089, 64090, 
    64091, 64092, 64093, 64094, 64095, 64096, 64097, 64098, 64099, 64100, 
    64101, 64102, 64103, 64104, 64105, 64106, 64107, 64108, 64109, 64110, 
    64111, 64112, 64113, 64114, 64115, 64116, 64117, 64118, 64119, 64120, 
    64121, 64122, 64123, 64124, 64125, 64126, 64127, 64128, 64129, 64130, 
    64131, 64132, 64133, 64134, 64135, 64136, 64137, 64138, 64139, 64140, 
    64141, 64142, 64143, 64144, 64145, 64146, 64147, 64148, 64149, 64150, 
    64151, 64152, 64153, 64154, 64155, 64156, 64157, 64158, 64159, 64160, 
    64161, 64162, 64163, 64164, 64165, 64166, 64167, 64168, 64169, 64170, 
    64171, 64172, 64173, 64174, 64175, 64176, 64177, 64178, 64179, 64180, 
    64181, 64182, 64183, 64184, 64185, 64186, 64187, 64188, 64189, 64190, 
    64191, 64192, 64193, 64194, 64195, 64196, 64197, 64198, 64199, 64200, 
    64201, 64202, 64203, 64204, 64205, 64206, 64207, 64208, 64209, 64210, 
    64211, 64212, 64213, 64214, 64215, 64216, 64217, 64218, 64219, 64220, 
    64221, 64222, 64223, 64224, 64225, 64226, 64227, 64228, 64229, 64230, 
    64231, 64232, 64233, 64234, 64235, 64236, 64237, 64238, 64239, 64240, 
    64241, 64242, 64243, 64244, 64245, 64246, 64247, 64248, 64249, 64250, 
    64251, 64252, 64253, 64254, 64255, 64256, 64257, 64258, 64259, 64260, 
    64261, 64262, 64263, 64264, 64265, 64266, 64267, 64268, 64269, 64270, 
    64271, 64272, 64273, 64274, 64275, 64276, 64277, 64278, 64279, 64280, 
    64281, 64282, 64283, 64284, 64285, 64286, 64287, 64288, 64289, 64290, 
    64291, 64292, 64293, 64294, 64295, 64296, 64297, 64298, 64299, 64300, 
    64301, 64302, 64303, 64304, 64305, 64306, 64307, 64308, 64309, 64310, 
    64311, 64312, 64313, 64314, 64315, 64316, 64317, 64318, 64319, 64320, 
    64321, 64322, 64323, 64324, 64325, 64326, 64327, 64328, 64329, 64330, 
    64331, 64332, 64333, 64334, 64335, 64336, 64337, 64338, 64339, 64340, 
    64341, 64342, 64343, 64344, 64345, 64346, 64347, 64348, 64349, 64350, 
    64351, 64352, 64353, 64354, 64355, 64356, 64357, 64358, 64359, 64360, 
    64361, 64362, 64363, 64364, 64365, 64366, 64367, 64368, 64369, 64370, 
    64371, 64372, 64373, 64374, 64375, 64376, 64377, 64378, 64379, 64380, 
    64381, 64382, 64383, 64384, 64385, 64386, 64387, 64388, 64389, 64390, 
    64391, 64392, 64393, 64394, 64395, 64396, 64397, 64398, 64399, 64400, 
    64401, 64402, 64403, 64404, 64405, 64406, 64407, 64408, 64409, 64410, 
    64411, 64412, 64413, 64414, 64415, 64416, 64417, 64418, 64419, 64420, 
    64421, 64422, 64423, 64424, 64425, 64426, 64427, 64428, 64429, 64430, 
    64431, 64432, 64433, 64434, 64435, 64436, 64437, 64438, 64439, 64440, 
    64441, 64442, 64443, 64444, 64445, 64446, 64447, 64448, 64449, 64450, 
    64451, 64452, 64453, 64454, 64455, 64456, 64457, 64458, 64459, 64460, 
    64461, 64462, 64463, 64464, 64465, 64466, 64467, 64468, 64469, 64470, 
    64471, 64472, 64473, 64474, 64475, 64476, 64477, 64478, 64479, 64480, 
    64481, 64482, 64483, 64484, 64485, 64486, 64487, 64488, 64489, 64490, 
    64491, 64492, 64493, 64494, 64495, 64496, 64497, 64498, 64499, 64500, 
    64501, 64502, 64503, 64504, 64505, 64506, 64507, 64508, 64509, 64510, 
    64511, 64512, 64513, 64514, 64515, 64516, 64517, 64518, 64519, 64520, 
    64521, 64522, 64523, 64524, 64525, 64526, 64527, 64528, 64529, 64530, 
    64531, 64532, 64533, 64534, 64535, 64536, 64537, 64538, 64539, 64540, 
    64541, 64542, 64543, 64544, 64545, 64546, 64547, 64548, 64549, 64550, 
    64551, 64552, 64553, 64554, 64555, 64556, 64557, 64558, 64559, 64560, 
    64561, 64562, 64563, 64564, 64565, 64566, 64567, 64568, 64569, 64570, 
    64571, 64572, 64573, 64574, 64575, 64576, 64577, 64578, 64579, 64580, 
    64581, 64582, 64583, 64584, 64585, 64586, 64587, 64588, 64589, 64590, 
    64591, 64592, 64593, 64594, 64595, 64596, 64597, 64598, 64599, 64600, 
    64601, 64602, 64603, 64604, 64605, 64606, 64607, 64608, 64609, 64610, 
    64611, 64612, 64613, 64614, 64615, 64616, 64617, 64618, 64619, 64620, 
    64621, 64622, 64623, 64624, 64625, 64626, 64627, 64628, 64629, 64630, 
    64631, 64632, 64633, 64634, 64635, 64636, 64637, 64638, 64639, 64640, 
    64641, 64642, 64643, 64644, 64645, 64646, 64647, 64648, 64649, 64650, 
    64651, 64652, 64653, 64654, 64655, 64656, 64657, 64658, 64659, 64660, 
    64661, 64662, 64663, 64664, 64665, 64666, 64667, 64668, 64669, 64670, 
    64671, 64672, 64673, 64674, 64675, 64676, 64677, 64678, 64679, 64680, 
    64681, 64682, 64683, 64684, 64685, 64686, 64687, 64688, 64689, 64690, 
    64691, 64692, 64693, 64694, 64695, 64696, 64697, 64698, 64699, 64700, 
    64701, 64702, 64703, 64704, 64705, 64706, 64707, 64708, 64709, 64710, 
    64711, 64712, 64713, 64714, 64715, 64716, 64717, 64718, 64719, 64720, 
    64721, 64722, 64723, 64724, 64725, 64726, 64727, 64728, 64729, 64730, 
    64731, 64732, 64733, 64734, 64735, 64736, 64737, 64738, 64739, 64740, 
    64741, 64742, 64743, 64744, 64745, 64746, 64747, 64748, 64749, 64750, 
    64751, 64752, 64753, 64754, 64755, 64756, 64757, 64758, 64759, 64760, 
    64761, 64762, 64763, 64764, 64765, 64766, 64767, 64768, 64769, 64770, 
    64771, 64772, 64773, 64774, 64775, 64776, 64777, 64778, 64779, 64780, 
    64781, 64782, 64783, 64784, 64785, 64786, 64787, 64788, 64789, 64790, 
    64791, 64792, 64793, 64794, 64795, 64796, 64797, 64798, 64799, 64800, 
    64801, 64802, 64803, 64804, 64805, 64806, 64807, 64808, 64809, 64810, 
    64811, 64812, 64813, 64814, 64815, 64816, 64817, 64818, 64819, 64820, 
    64821, 64822, 64823, 64824, 64825, 64826, 64827, 64828, 64829, 64830, 
    64831, 64832, 64833, 64834, 64835, 64836, 64837, 64838, 64839, 64840, 
    64841, 64842, 64843, 64844, 64845, 64846, 64847, 64848, 64849, 64850, 
    64851, 64852, 64853, 64854, 64855, 64856, 64857, 64858, 64859, 64860, 
    64861, 64862, 64863, 64864, 64865, 64866, 64867, 64868, 64869, 64870, 
    64871, 64872, 64873, 64874, 64875, 64876, 64877, 64878, 64879, 64880, 
    64881, 64882, 64883, 64884, 64885, 64886, 64887, 64888, 64889, 64890, 
    64891, 64892, 64893, 64894, 64895, 64896, 64897, 64898, 64899, 64900, 
    64901, 64902, 64903, 64904, 64905, 64906, 64907, 64908, 64909, 64910, 
    64911, 64912, 64913, 64914, 64915, 64916, 64917, 64918, 64919, 64920, 
    64921, 64922, 64923, 64924, 64925, 64926, 64927, 64928, 64929, 64930, 
    64931, 64932, 64933, 64934, 64935, 64936, 64937, 64938, 64939, 64940, 
    64941, 64942, 64943, 64944, 64945, 64946, 64947, 64948, 64949, 64950, 
    64951, 64952, 64953, 64954, 64955, 64956, 64957, 64958, 64959, 64960, 
    64961, 64962, 64963, 64964, 64965, 64966, 64967, 64968, 64969, 64970, 
    64971, 64972, 64973, 64974, 64975, 64976, 64977, 64978, 64979, 64980, 
    64981, 64982, 64983, 64984, 64985, 64986, 64987, 64988, 64989, 64990, 
    64991, 64992, 64993, 64994, 64995, 64996, 64997, 64998, 64999, 65000, 
    65001, 65002, 65003, 65004, 65005, 65006, 65007, 65008, 65009, 65010, 
    65011, 65012, 65013, 65014, 65015, 65016, 65017, 65018, 65019, 65020, 
    65021, 65022, 65023, 65024, 65025, 65026, 65027, 65028, 65029, 65030, 
    65031, 65032, 65033, 65034, 65035, 65036, 65037, 65038, 65039, 65040, 
    65041, 65042, 65043, 65044, 65045, 65046, 65047, 65048, 65049, 65050, 
    65051, 65052, 65053, 65054, 65055, 65056, 65057, 65058, 65059, 65060, 
    65061, 65062, 65063, 65064, 65065, 65066, 65067, 65068, 65069, 65070, 
    65071, 65072, 65073, 65074, 65075, 65076, 65077, 65078, 65079, 65080, 
    65081, 65082, 65083, 65084, 65085, 65086, 65087, 65088, 65089, 65090, 
    65091, 65092, 65093, 65094, 65095, 65096, 65097, 65098, 65099, 65100, 
    65101, 65102, 65103, 65104, 65105, 65106, 65107, 65108, 65109, 65110, 
    65111, 65112, 65113, 65114, 65115, 65116, 65117, 65118, 65119, 65120, 
    65121, 65122, 65123, 65124, 65125, 65126, 65127, 65128, 65129, 65130, 
    65131, 65132, 65133, 65134, 65135, 65136, 65137, 65138, 65139, 65140, 
    65141, 65142, 65143, 65144, 65145, 65146, 65147, 65148, 65149, 65150, 
    65151, 65152, 65153, 65154, 65155, 65156, 65157, 65158, 65159, 65160, 
    65161, 65162, 65163, 65164, 65165, 65166, 65167, 65168, 65169, 65170, 
    65171, 65172, 65173, 65174, 65175, 65176, 65177, 65178, 65179, 65180, 
    65181, 65182, 65183, 65184, 65185, 65186, 65187, 65188, 65189, 65190, 
    65191, 65192, 65193, 65194, 65195, 65196, 65197, 65198, 65199, 65200, 
    65201, 65202, 65203, 65204, 65205, 65206, 65207, 65208, 65209, 65210, 
    65211, 65212, 65213, 65214, 65215, 65216, 65217, 65218, 65219, 65220, 
    65221, 65222, 65223, 65224, 65225, 65226, 65227, 65228, 65229, 65230, 
    65231, 65232, 65233, 65234, 65235, 65236, 65237, 65238, 65239, 65240, 
    65241, 65242, 65243, 65244, 65245, 65246, 65247, 65248, 65249, 65250, 
    65251, 65252, 65253, 65254, 65255, 65256, 65257, 65258, 65259, 65260, 
    65261, 65262, 65263, 65264, 65265, 65266, 65267, 65268, 65269, 65270, 
    65271, 65272, 65273, 65274, 65275, 65276, 65277, 65278, 65279, 65280, 
    65281, 65282, 65283, 65284, 65285, 65286, 65287, 65288, 65289, 65290, 
    65291, 65292, 65293, 65294, 65295, 65296, 65297, 65298, 65299, 65300, 
    65301, 65302, 65303, 65304, 65305, 65306, 65307, 65308, 65309, 65310, 
    65311, 65312, 65313, 65314, 65315, 65316, 65317, 65318, 65319, 65320, 
    65321, 65322, 65323, 65324, 65325, 65326, 65327, 65328, 65329, 65330, 
    65331, 65332, 65333, 65334, 65335, 65336, 65337, 65338, 65339, 65340, 
    65341, 65342, 65343, 65344, 65345, 65346, 65347, 65348, 65349, 65350, 
    65351, 65352, 65353, 65354, 65355, 65356, 65357, 65358, 65359, 65360, 
    65361, 65362, 65363, 65364, 65365, 65366, 65367, 65368, 65369, 65370, 
    65371, 65372, 65373, 65374, 65375, 65376, 65377, 65378, 65379, 65380, 
    65381, 65382, 65383, 65384, 65385, 65386, 65387, 65388, 65389, 65390, 
    65391, 65392, 65393, 65394, 65395, 65396, 65397, 65398, 65399, 65400, 
    65401, 65402, 65403, 65404, 65405, 65406, 65407, 65408, 65409, 65410, 
    65411, 65412, 65413, 65414, 65415, 65416, 65417, 65418, 65419, 65420, 
    65421, 65422, 65423, 65424, 65425, 65426, 65427, 65428, 65429, 65430, 
    65431, 65432, 65433, 65434, 65435, 65436, 65437, 65438, 65439, 65440, 
    65441, 65442, 65443, 65444, 65445, 65446, 65447, 65448, 65449, 65450, 
    65451, 65452, 65453, 65454, 65455, 65456, 65457, 65458, 65459, 65460, 
    65461, 65462, 65463, 65464, 65465, 65466, 65467, 65468, 65469, 65470, 
    65471, 65472, 65473, 65474, 65475, 65476, 65477, 65478, 65479, 65480, 
    65481, 65482, 65483, 65484, 65485, 65486, 65487, 65488, 65489, 65490, 
    65491, 65492, 65493, 65494, 65495, 65496, 65497, 65498, 65499, 65500, 
    65501, 65502, 65503, 65504, 65505, 65506, 65507, 65508, 65509, 65510, 
    65511, 65512, 65513, 65514, 65515, 65516, 65517, 65518, 65519, 65520, 
    65521, 65522, 65523, 65524, 65525, 65526, 65527, 65528, 65529, 65530, 
    65531, 65532, 65533, 65534, 65535, 65536, 65537, 65538, 65539, 65540, 
    65541, 65542, 65543, 65544, 65545, 65546, 65547, 65548, 65549, 65550, 
    65551, 65552, 65553, 65554, 65555, 65556, 65557, 65558, 65559, 65560, 
    65561, 65562, 65563, 65564, 65565, 65566, 65567, 65568, 65569, 65570, 
    65571, 65572, 65573, 65574, 65575, 65576, 65577, 65578, 65579, 65580, 
    65581, 65582, 65583, 65584, 65585, 65586, 65587, 65588, 65589, 65590, 
    65591, 65592, 65593, 65594, 65595, 65596, 65597, 65598, 65599, 65600, 
    65601, 65602, 65603, 65604, 65605, 65606, 65607, 65608, 65609, 65610, 
    65611, 65612, 65613, 65614, 65615, 65616, 65617, 65618, 65619, 65620, 
    65621, 65622, 65623, 65624, 65625, 65626, 65627, 65628, 65629, 65630, 
    65631, 65632, 65633, 65634, 65635, 65636, 65637, 65638, 65639, 65640, 
    65641, 65642, 65643, 65644, 65645, 65646, 65647, 65648, 65649, 65650, 
    65651, 65652, 65653, 65654, 65655, 65656, 65657, 65658, 65659, 65660, 
    65661, 65662, 65663, 65664, 65665, 65666, 65667, 65668, 65669, 65670, 
    65671, 65672, 65673, 65674, 65675, 65676, 65677, 65678, 65679, 65680, 
    65681, 65682, 65683, 65684, 65685, 65686, 65687, 65688, 65689, 65690, 
    65691, 65692, 65693, 65694, 65695, 65696, 65697, 65698, 65699, 65700, 
    65701, 65702, 65703, 65704, 65705, 65706, 65707, 65708, 65709, 65710, 
    65711, 65712, 65713, 65714, 65715, 65716, 65717, 65718, 65719, 65720, 
    65721, 65722, 65723, 65724, 65725, 65726, 65727, 65728, 65729, 65730, 
    65731, 65732, 65733, 65734, 65735, 65736, 65737, 65738, 65739, 65740, 
    65741, 65742, 65743, 65744, 65745, 65746, 65747, 65748, 65749, 65750, 
    65751, 65752, 65753, 65754, 65755, 65756, 65757, 65758, 65759, 65760, 
    65761, 65762, 65763, 65764, 65765, 65766, 65767, 65768, 65769, 65770, 
    65771, 65772, 65773, 65774, 65775, 65776, 65777, 65778, 65779, 65780, 
    65781, 65782, 65783, 65784, 65785, 65786, 65787, 65788, 65789, 65790, 
    65791, 65792, 65793, 65794, 65795, 65796, 65797, 65798, 65799, 65800, 
    65801, 65802, 65803, 65804, 65805, 65806, 65807, 65808, 65809, 65810, 
    65811, 65812, 65813, 65814, 65815, 65816, 65817, 65818, 65819, 65820, 
    65821, 65822, 65823, 65824, 65825, 65826, 65827, 65828, 65829, 65830, 
    65831, 65832, 65833, 65834, 65835, 65836, 65837, 65838, 65839, 65840, 
    65841, 65842, 65843, 65844, 65845, 65846, 65847, 65848, 65849, 65850, 
    65851, 65852, 65853, 65854, 65855, 65856, 65857, 65858, 65859, 65860, 
    65861, 65862, 65863, 65864, 65865, 65866, 65867, 65868, 65869, 65870, 
    65871, 65872, 65873, 65874, 65875, 65876, 65877, 65878, 65879, 65880, 
    65881, 65882, 65883, 65884, 65885, 65886, 65887, 65888, 65889, 65890, 
    65891, 65892, 65893, 65894, 65895, 65896, 65897, 65898, 65899, 65900, 
    65901, 65902, 65903, 65904, 65905, 65906, 65907, 65908, 65909, 65910, 
    65911, 65912, 65913, 65914, 65915, 65916, 65917, 65918, 65919, 65920, 
    65921, 65922, 65923, 65924, 65925, 65926, 65927, 65928, 65929, 65930, 
    65931, 65932, 65933, 65934, 65935, 65936, 65937, 65938, 65939, 65940, 
    65941, 65942, 65943, 65944, 65945, 65946, 65947, 65948, 65949, 65950, 
    65951, 65952, 65953, 65954, 65955, 65956, 65957, 65958, 65959, 65960, 
    65961, 65962, 65963, 65964, 65965, 65966, 65967, 65968, 65969, 65970, 
    65971, 65972, 65973, 65974, 65975, 65976, 65977, 65978, 65979, 65980, 
    65981, 65982, 65983, 65984, 65985, 65986, 65987, 65988, 65989, 65990, 
    65991, 65992, 65993, 65994, 65995, 65996, 65997, 65998, 65999, 66000, 
    66001, 66002, 66003, 66004, 66005, 66006, 66007, 66008, 66009, 66010, 
    66011, 66012, 66013, 66014, 66015, 66016, 66017, 66018, 66019, 66020, 
    66021, 66022, 66023, 66024, 66025, 66026, 66027, 66028, 66029, 66030, 
    66031, 66032, 66033, 66034, 66035, 66036, 66037, 66038, 66039, 66040, 
    66041, 66042, 66043, 66044, 66045, 66046, 66047, 66048, 66049, 66050, 
    66051, 66052, 66053, 66054, 66055, 66056, 66057, 66058, 66059, 66060, 
    66061, 66062, 66063, 66064, 66065, 66066, 66067, 66068, 66069, 66070, 
    66071, 66072, 66073, 66074, 66075, 66076, 66077, 66078, 66079, 66080, 
    66081, 66082, 66083, 66084, 66085, 66086, 66087, 66088, 66089, 66090, 
    66091, 66092, 66093, 66094, 66095, 66096, 66097, 66098, 66099, 66100, 
    66101, 66102, 66103, 66104, 66105, 66106, 66107, 66108, 66109, 66110, 
    66111, 66112, 66113, 66114, 66115, 66116, 66117, 66118, 66119, 66120, 
    66121, 66122, 66123, 66124, 66125, 66126, 66127, 66128, 66129, 66130, 
    66131, 66132, 66133, 66134, 66135, 66136, 66137, 66138, 66139, 66140, 
    66141, 66142, 66143, 66144, 66145, 66146, 66147, 66148, 66149, 66150, 
    66151, 66152, 66153, 66154, 66155, 66156, 66157, 66158, 66159, 66160, 
    66161, 66162, 66163, 66164, 66165, 66166, 66167, 66168, 66169, 66170, 
    66171, 66172, 66173, 66174, 66175, 66176, 66177, 66178, 66179, 66180, 
    66181, 66182, 66183, 66184, 66185, 66186, 66187, 66188, 66189, 66190, 
    66191, 66192, 66193, 66194, 66195, 66196, 66197, 66198, 66199, 66200, 
    66201, 66202, 66203, 66204, 66205, 66206, 66207, 66208, 66209, 66210, 
    66211, 66212, 66213, 66214, 66215, 66216, 66217, 66218, 66219, 66220, 
    66221, 66222, 66223, 66224, 66225, 66226, 66227, 66228, 66229, 66230, 
    66231, 66232, 66233, 66234, 66235, 66236, 66237, 66238, 66239, 66240, 
    66241, 66242, 66243, 66244, 66245, 66246, 66247, 66248, 66249, 66250, 
    66251, 66252, 66253, 66254, 66255, 66256, 66257, 66258, 66259, 66260, 
    66261, 66262, 66263, 66264, 66265, 66266, 66267, 66268, 66269, 66270, 
    66271, 66272, 66273, 66274, 66275, 66276, 66277, 66278, 66279, 66280, 
    66281, 66282, 66283, 66284, 66285, 66286, 66287, 66288, 66289, 66290, 
    66291, 66292, 66293, 66294, 66295, 66296, 66297, 66298, 66299, 66300, 
    66301, 66302, 66303, 66304, 66305, 66306, 66307, 66308, 66309, 66310, 
    66311, 66312, 66313, 66314, 66315, 66316, 66317, 66318, 66319, 66320, 
    66321, 66322, 66323, 66324, 66325, 66326, 66327, 66328, 66329, 66330, 
    66331, 66332, 66333, 66334, 66335, 66336, 66337, 66338, 66339, 66340, 
    66341, 66342, 66343, 66344, 66345, 66346, 66347, 66348, 66349, 66350, 
    66351, 66352, 66353, 66354, 66355, 66356, 66357, 66358, 66359, 66360, 
    66361, 66362, 66363, 66364, 66365, 66366, 66367, 66368, 66369, 66370, 
    66371, 66372, 66373, 66374, 66375, 66376, 66377, 66378, 66379, 66380, 
    66381, 66382, 66383, 66384, 66385, 66386, 66387, 66388, 66389, 66390, 
    66391, 66392, 66393, 66394, 66395, 66396, 66397, 66398, 66399, 66400, 
    66401, 66402, 66403, 66404, 66405, 66406, 66407, 66408, 66409, 66410, 
    66411, 66412, 66413, 66414, 66415, 66416, 66417, 66418, 66419, 66420, 
    66421, 66422, 66423, 66424, 66425, 66426, 66427, 66428, 66429, 66430, 
    66431, 66432, 66433, 66434, 66435, 66436, 66437, 66438, 66439, 66440, 
    66441, 66442, 66443, 66444, 66445, 66446, 66447, 66448, 66449, 66450, 
    66451, 66452, 66453, 66454, 66455, 66456, 66457, 66458, 66459, 66460, 
    66461, 66462, 66463, 66464, 66465, 66466, 66467, 66468, 66469, 66470, 
    66471, 66472, 66473, 66474, 66475, 66476, 66477, 66478, 66479, 66480, 
    66481, 66482, 66483, 66484, 66485, 66486, 66487, 66488, 66489, 66490, 
    66491, 66492, 66493, 66494, 66495, 66496, 66497, 66498, 66499, 66500, 
    66501, 66502, 66503, 66504, 66505, 66506, 66507, 66508, 66509, 66510, 
    66511, 66512, 66513, 66514, 66515, 66516, 66517, 66518, 66519, 66520, 
    66521, 66522, 66523, 66524, 66525, 66526, 66527, 66528, 66529, 66530, 
    66531, 66532, 66533, 66534, 66535, 66536, 66537, 66538, 66539, 66540, 
    66541, 66542, 66543, 66544, 66545, 66546, 66547, 66548, 66549, 66550, 
    66551, 66552, 66553, 66554, 66555, 66556, 66557, 66558, 66559, 66560, 
    66561, 66562, 66563, 66564, 66565, 66566, 66567, 66568, 66569, 66570, 
    66571, 66572, 66573, 66574, 66575, 66576, 66577, 66578, 66579, 66580, 
    66581, 66582, 66583, 66584, 66585, 66586, 66587, 66588, 66589, 66590, 
    66591, 66592, 66593, 66594, 66595, 66596, 66597, 66598, 66599, 66600, 
    66601, 66602, 66603, 66604, 66605, 66606, 66607, 66608, 66609, 66610, 
    66611, 66612, 66613, 66614, 66615, 66616, 66617, 66618, 66619, 66620, 
    66621, 66622, 66623, 66624, 66625, 66626, 66627, 66628, 66629, 66630, 
    66631, 66632, 66633, 66634, 66635, 66636, 66637, 66638, 66639, 66640, 
    66641, 66642, 66643, 66644, 66645, 66646, 66647, 66648, 66649, 66650, 
    66651, 66652, 66653, 66654, 66655, 66656, 66657, 66658, 66659, 66660, 
    66661, 66662, 66663, 66664, 66665, 66666, 66667, 66668, 66669, 66670, 
    66671, 66672, 66673, 66674, 66675, 66676, 66677, 66678, 66679, 66680, 
    66681, 66682, 66683, 66684, 66685, 66686, 66687, 66688, 66689, 66690, 
    66691, 66692, 66693, 66694, 66695, 66696, 66697, 66698, 66699, 66700, 
    66701, 66702, 66703, 66704, 66705, 66706, 66707, 66708, 66709, 66710, 
    66711, 66712, 66713, 66714, 66715, 66716, 66717, 66718, 66719, 66720, 
    66721, 66722, 66723, 66724, 66725, 66726, 66727, 66728, 66729, 66730, 
    66731, 66732, 66733, 66734, 66735, 66736, 66737, 66738, 66739, 66740, 
    66741, 66742, 66743, 66744, 66745, 66746, 66747, 66748, 66749, 66750, 
    66751, 66752, 66753, 66754, 66755, 66756, 66757, 66758, 66759, 66760, 
    66761, 66762, 66763, 66764, 66765, 66766, 66767, 66768, 66769, 66770, 
    66771, 66772, 66773, 66774, 66775, 66776, 66777, 66778, 66779, 66780, 
    66781, 66782, 66783, 66784, 66785, 66786, 66787, 66788, 66789, 66790, 
    66791, 66792, 66793, 66794, 66795, 66796, 66797, 66798, 66799, 66800, 
    66801, 66802, 66803, 66804, 66805, 66806, 66807, 66808, 66809, 66810, 
    66811, 66812, 66813, 66814, 66815, 66816, 66817, 66818, 66819, 66820, 
    66821, 66822, 66823, 66824, 66825, 66826, 66827, 66828, 66829, 66830, 
    66831, 66832, 66833, 66834, 66835, 66836, 66837, 66838, 66839, 66840, 
    66841, 66842, 66843, 66844, 66845, 66846, 66847, 66848, 66849, 66850, 
    66851, 66852, 66853, 66854, 66855, 66856, 66857, 66858, 66859, 66860, 
    66861, 66862, 66863, 66864, 66865, 66866, 66867, 66868, 66869, 66870, 
    66871, 66872, 66873, 66874, 66875, 66876, 66877, 66878, 66879, 66880, 
    66881, 66882, 66883, 66884, 66885, 66886, 66887, 66888, 66889, 66890, 
    66891, 66892, 66893, 66894, 66895, 66896, 66897, 66898, 66899, 66900, 
    66901, 66902, 66903, 66904, 66905, 66906, 66907, 66908, 66909, 66910, 
    66911, 66912, 66913, 66914, 66915, 66916, 66917, 66918, 66919, 66920, 
    66921, 66922, 66923, 66924, 66925, 66926, 66927, 66928, 66929, 66930, 
    66931, 66932, 66933, 66934, 66935, 66936, 66937, 66938, 66939, 66940, 
    66941, 66942, 66943, 66944, 66945, 66946, 66947, 66948, 66949, 66950, 
    66951, 66952, 66953, 66954, 66955, 66956, 66957, 66958, 66959, 66960, 
    66961, 66962, 66963, 66964, 66965, 66966, 66967, 66968, 66969, 66970, 
    66971, 66972, 66973, 66974, 66975, 66976, 66977, 66978, 66979, 66980, 
    66981, 66982, 66983, 66984, 66985, 66986, 66987, 66988, 66989, 66990, 
    66991, 66992, 66993, 66994, 66995, 66996, 66997, 66998, 66999, 67000, 
    67001, 67002, 67003, 67004, 67005, 67006, 67007, 67008, 67009, 67010, 
    67011, 67012, 67013, 67014, 67015, 67016, 67017, 67018, 67019, 67020, 
    67021, 67022, 67023, 67024, 67025, 67026, 67027, 67028, 67029, 67030, 
    67031, 67032, 67033, 67034, 67035, 67036, 67037, 67038, 67039, 67040, 
    67041, 67042, 67043, 67044, 67045, 67046, 67047, 67048, 67049, 67050, 
    67051, 67052, 67053, 67054, 67055, 67056, 67057, 67058, 67059, 67060, 
    67061, 67062, 67063, 67064, 67065, 67066, 67067, 67068, 67069, 67070, 
    67071, 67072, 67073, 67074, 67075, 67076, 67077, 67078, 67079, 67080, 
    67081, 67082, 67083, 67084, 67085, 67086, 67087, 67088, 67089, 67090, 
    67091, 67092, 67093, 67094, 67095, 67096, 67097, 67098, 67099, 67100, 
    67101, 67102, 67103, 67104, 67105, 67106, 67107, 67108, 67109, 67110, 
    67111, 67112, 67113, 67114, 67115, 67116, 67117, 67118, 67119, 67120, 
    67121, 67122, 67123, 67124, 67125, 67126, 67127, 67128, 67129, 67130, 
    67131, 67132, 67133, 67134, 67135, 67136, 67137, 67138, 67139, 67140, 
    67141, 67142, 67143, 67144, 67145, 67146, 67147, 67148, 67149, 67150, 
    67151, 67152, 67153, 67154, 67155, 67156, 67157, 67158, 67159, 67160, 
    67161, 67162, 67163, 67164, 67165, 67166, 67167, 67168, 67169, 67170, 
    67171, 67172, 67173, 67174, 67175, 67176, 67177, 67178, 67179, 67180, 
    67181, 67182, 67183, 67184, 67185, 67186, 67187, 67188, 67189, 67190, 
    67191, 67192, 67193, 67194, 67195, 67196, 67197, 67198, 67199, 67200, 
    67201, 67202, 67203, 67204, 67205, 67206, 67207, 67208, 67209, 67210, 
    67211, 67212, 67213, 67214, 67215, 67216, 67217, 67218, 67219, 67220, 
    67221, 67222, 67223, 67224, 67225, 67226, 67227, 67228, 67229, 67230, 
    67231, 67232, 67233, 67234, 67235, 67236, 67237, 67238, 67239, 67240, 
    67241, 67242, 67243, 67244, 67245, 67246, 67247, 67248, 67249, 67250, 
    67251, 67252, 67253, 67254, 67255, 67256, 67257, 67258, 67259, 67260, 
    67261, 67262, 67263, 67264, 67265, 67266, 67267, 67268, 67269, 67270, 
    67271, 67272, 67273, 67274, 67275, 67276, 67277, 67278, 67279, 67280, 
    67281, 67282, 67283, 67284, 67285, 67286, 67287, 67288, 67289, 67290, 
    67291, 67292, 67293, 67294, 67295, 67296, 67297, 67298, 67299, 67300, 
    67301, 67302, 67303, 67304, 67305, 67306, 67307, 67308, 67309, 67310, 
    67311, 67312, 67313, 67314, 67315, 67316, 67317, 67318, 67319, 67320, 
    67321, 67322, 67323, 67324, 67325, 67326, 67327, 67328, 67329, 67330, 
    67331, 67332, 67333, 67334, 67335, 67336, 67337, 67338, 67339, 67340, 
    67341, 67342, 67343, 67344, 67345, 67346, 67347, 67348, 67349, 67350, 
    67351, 67352, 67353, 67354, 67355, 67356, 67357, 67358, 67359, 67360, 
    67361, 67362, 67363, 67364, 67365, 67366, 67367, 67368, 67369, 67370, 
    67371, 67372, 67373, 67374, 67375, 67376, 67377, 67378, 67379, 67380, 
    67381, 67382, 67383, 67384, 67385, 67386, 67387, 67388, 67389, 67390, 
    67391, 67392, 67393, 67394, 67395, 67396, 67397, 67398, 67399, 67400, 
    67401, 67402, 67403, 67404, 67405, 67406, 67407, 67408, 67409, 67410, 
    67411, 67412, 67413, 67414, 67415, 67416, 67417, 67418, 67419, 67420, 
    67421, 67422, 67423, 67424, 67425, 67426, 67427, 67428, 67429, 67430, 
    67431, 67432, 67433, 67434, 67435, 67436, 67437, 67438, 67439, 67440, 
    67441, 67442, 67443, 67444, 67445, 67446, 67447, 67448, 67449, 67450, 
    67451, 67452, 67453, 67454, 67455, 67456, 67457, 67458, 67459, 67460, 
    67461, 67462, 67463, 67464, 67465, 67466, 67467, 67468, 67469, 67470, 
    67471, 67472, 67473, 67474, 67475, 67476, 67477, 67478, 67479, 67480, 
    67481, 67482, 67483, 67484, 67485, 67486, 67487, 67488, 67489, 67490, 
    67491, 67492, 67493, 67494, 67495, 67496, 67497, 67498, 67499, 67500, 
    67501, 67502, 67503, 67504, 67505, 67506, 67507, 67508, 67509, 67510, 
    67511, 67512, 67513, 67514, 67515, 67516, 67517, 67518, 67519, 67520, 
    67521, 67522, 67523, 67524, 67525, 67526, 67527, 67528, 67529, 67530, 
    67531, 67532, 67533, 67534, 67535, 67536, 67537, 67538, 67539, 67540, 
    67541, 67542, 67543, 67544, 67545, 67546, 67547, 67548, 67549, 67550, 
    67551, 67552, 67553, 67554, 67555, 67556, 67557, 67558, 67559, 67560, 
    67561, 67562, 67563, 67564, 67565, 67566, 67567, 67568, 67569, 67570, 
    67571, 67572, 67573, 67574, 67575, 67576, 67577, 67578, 67579, 67580, 
    67581, 67582, 67583, 67584, 67585, 67586, 67587, 67588, 67589, 67590, 
    67591, 67592, 67593, 67594, 67595, 67596, 67597, 67598, 67599, 67600, 
    67601, 67602, 67603, 67604, 67605, 67606, 67607, 67608, 67609, 67610, 
    67611, 67612, 67613, 67614, 67615, 67616, 67617, 67618, 67619, 67620, 
    67621, 67622, 67623, 67624, 67625, 67626, 67627, 67628, 67629, 67630, 
    67631, 67632, 67633, 67634, 67635, 67636, 67637, 67638, 67639, 67640, 
    67641, 67642, 67643, 67644, 67645, 67646, 67647, 67648, 67649, 67650, 
    67651, 67652, 67653, 67654, 67655, 67656, 67657, 67658, 67659, 67660, 
    67661, 67662, 67663, 67664, 67665, 67666, 67667, 67668, 67669, 67670, 
    67671, 67672, 67673, 67674, 67675, 67676, 67677, 67678, 67679, 67680, 
    67681, 67682, 67683, 67684, 67685, 67686, 67687, 67688, 67689, 67690, 
    67691, 67692, 67693, 67694, 67695, 67696, 67697, 67698, 67699, 67700, 
    67701, 67702, 67703, 67704, 67705, 67706, 67707, 67708, 67709, 67710, 
    67711, 67712, 67713, 67714, 67715, 67716, 67717, 67718, 67719, 67720, 
    67721, 67722, 67723, 67724, 67725, 67726, 67727, 67728, 67729, 67730, 
    67731, 67732, 67733, 67734, 67735, 67736, 67737, 67738, 67739, 67740, 
    67741, 67742, 67743, 67744, 67745, 67746, 67747, 67748, 67749, 67750, 
    67751, 67752, 67753, 67754, 67755, 67756, 67757, 67758, 67759, 67760, 
    67761, 67762, 67763, 67764, 67765, 67766, 67767, 67768, 67769, 67770, 
    67771, 67772, 67773, 67774, 67775, 67776, 67777, 67778, 67779, 67780, 
    67781, 67782, 67783, 67784, 67785, 67786, 67787, 67788, 67789, 67790, 
    67791, 67792, 67793, 67794, 67795, 67796, 67797, 67798, 67799, 67800, 
    67801, 67802, 67803, 67804, 67805, 67806, 67807, 67808, 67809, 67810, 
    67811, 67812, 67813, 67814, 67815, 67816, 67817, 67818, 67819, 67820, 
    67821, 67822, 67823, 67824, 67825, 67826, 67827, 67828, 67829, 67830, 
    67831, 67832, 67833, 67834, 67835, 67836, 67837, 67838, 67839, 67840, 
    67841, 67842, 67843, 67844, 67845, 67846, 67847, 67848, 67849, 67850, 
    67851, 67852, 67853, 67854, 67855, 67856, 67857, 67858, 67859, 67860, 
    67861, 67862, 67863, 67864, 67865, 67866, 67867, 67868, 67869, 67870, 
    67871, 67872, 67873, 67874, 67875, 67876, 67877, 67878, 67879, 67880, 
    67881, 67882, 67883, 67884, 67885, 67886, 67887, 67888, 67889, 67890, 
    67891, 67892, 67893, 67894, 67895, 67896, 67897, 67898, 67899, 67900, 
    67901, 67902, 67903, 67904, 67905, 67906, 67907, 67908, 67909, 67910, 
    67911, 67912, 67913, 67914, 67915, 67916, 67917, 67918, 67919, 67920, 
    67921, 67922, 67923, 67924, 67925, 67926, 67927, 67928, 67929, 67930, 
    67931, 67932, 67933, 67934, 67935, 67936, 67937, 67938, 67939, 67940, 
    67941, 67942, 67943, 67944, 67945, 67946, 67947, 67948, 67949, 67950, 
    67951, 67952, 67953, 67954, 67955, 67956, 67957, 67958, 67959, 67960, 
    67961, 67962, 67963, 67964, 67965, 67966, 67967, 67968, 67969, 67970, 
    67971, 67972, 67973, 67974, 67975, 67976, 67977, 67978, 67979, 67980, 
    67981, 67982, 67983, 67984, 67985, 67986, 67987, 67988, 67989, 67990, 
    67991, 67992, 67993, 67994, 67995, 67996, 67997, 67998, 67999, 68000, 
    68001, 68002, 68003, 68004, 68005, 68006, 68007, 68008, 68009, 68010, 
    68011, 68012, 68013, 68014, 68015, 68016, 68017, 68018, 68019, 68020, 
    68021, 68022, 68023, 68024, 68025, 68026, 68027, 68028, 68029, 68030, 
    68031, 68032, 68033, 68034, 68035, 68036, 68037, 68038, 68039, 68040, 
    68041, 68042, 68043, 68044, 68045, 68046, 68047, 68048, 68049, 68050, 
    68051, 68052, 68053, 68054, 68055, 68056, 68057, 68058, 68059, 68060, 
    68061, 68062, 68063, 68064, 68065, 68066, 68067, 68068, 68069, 68070, 
    68071, 68072, 68073, 68074, 68075, 68076, 68077, 68078, 68079, 68080, 
    68081, 68082, 68083, 68084, 68085, 68086, 68087, 68088, 68089, 68090, 
    68091, 68092, 68093, 68094, 68095, 68096, 68097, 68098, 68099, 68100, 
    68101, 68102, 68103, 68104, 68105, 68106, 68107, 68108, 68109, 68110, 
    68111, 68112, 68113, 68114, 68115, 68116, 68117, 68118, 68119, 68120, 
    68121, 68122, 68123, 68124, 68125, 68126, 68127, 68128, 68129, 68130, 
    68131, 68132, 68133, 68134, 68135, 68136, 68137, 68138, 68139, 68140, 
    68141, 68142, 68143, 68144, 68145, 68146, 68147, 68148, 68149, 68150, 
    68151, 68152, 68153, 68154, 68155, 68156, 68157, 68158, 68159, 68160, 
    68161, 68162, 68163, 68164, 68165, 68166, 68167, 68168, 68169, 68170, 
    68171, 68172, 68173, 68174, 68175, 68176, 68177, 68178, 68179, 68180, 
    68181, 68182, 68183, 68184, 68185, 68186, 68187, 68188, 68189, 68190, 
    68191, 68192, 68193, 68194, 68195, 68196, 68197, 68198, 68199, 68200, 
    68201, 68202, 68203, 68204, 68205, 68206, 68207, 68208, 68209, 68210, 
    68211, 68212, 68213, 68214, 68215, 68216, 68217, 68218, 68219, 68220, 
    68221, 68222, 68223, 68224, 68225, 68226, 68227, 68228, 68229, 68230, 
    68231, 68232, 68233, 68234, 68235, 68236, 68237, 68238, 68239, 68240, 
    68241, 68242, 68243, 68244, 68245, 68246, 68247, 68248, 68249, 68250, 
    68251, 68252, 68253, 68254, 68255, 68256, 68257, 68258, 68259, 68260, 
    68261, 68262, 68263, 68264, 68265, 68266, 68267, 68268, 68269, 68270, 
    68271, 68272, 68273, 68274, 68275, 68276, 68277, 68278, 68279, 68280, 
    68281, 68282, 68283, 68284, 68285, 68286, 68287, 68288, 68289, 68290, 
    68291, 68292, 68293, 68294, 68295, 68296, 68297, 68298, 68299, 68300, 
    68301, 68302, 68303, 68304, 68305, 68306, 68307, 68308, 68309, 68310, 
    68311, 68312, 68313, 68314, 68315, 68316, 68317, 68318, 68319, 68320, 
    68321, 68322, 68323, 68324, 68325, 68326, 68327, 68328, 68329, 68330, 
    68331, 68332, 68333, 68334, 68335, 68336, 68337, 68338, 68339, 68340, 
    68341, 68342, 68343, 68344, 68345, 68346, 68347, 68348, 68349, 68350, 
    68351, 68352, 68353, 68354, 68355, 68356, 68357, 68358, 68359, 68360, 
    68361, 68362, 68363, 68364, 68365, 68366, 68367, 68368, 68369, 68370, 
    68371, 68372, 68373, 68374, 68375, 68376, 68377, 68378, 68379, 68380, 
    68381, 68382, 68383, 68384, 68385, 68386, 68387, 68388, 68389, 68390, 
    68391, 68392, 68393, 68394, 68395, 68396, 68397, 68398, 68399, 68400, 
    68401, 68402, 68403, 68404, 68405, 68406, 68407, 68408, 68409, 68410, 
    68411, 68412, 68413, 68414, 68415, 68416, 68417, 68418, 68419, 68420, 
    68421, 68422, 68423, 68424, 68425, 68426, 68427, 68428, 68429, 68430, 
    68431, 68432, 68433, 68434, 68435, 68436, 68437, 68438, 68439, 68440, 
    68441, 68442, 68443, 68444, 68445, 68446, 68447, 68448, 68449, 68450, 
    68451, 68452, 68453, 68454, 68455, 68456, 68457, 68458, 68459, 68460, 
    68461, 68462, 68463, 68464, 68465, 68466, 68467, 68468, 68469, 68470, 
    68471, 68472, 68473, 68474, 68475, 68476, 68477, 68478, 68479, 68480, 
    68481, 68482, 68483, 68484, 68485, 68486, 68487, 68488, 68489, 68490, 
    68491, 68492, 68493, 68494, 68495, 68496, 68497, 68498, 68499, 68500, 
    68501, 68502, 68503, 68504, 68505, 68506, 68507, 68508, 68509, 68510, 
    68511, 68512, 68513, 68514, 68515, 68516, 68517, 68518, 68519, 68520, 
    68521, 68522, 68523, 68524, 68525, 68526, 68527, 68528, 68529, 68530, 
    68531, 68532, 68533, 68534, 68535, 68536, 68537, 68538, 68539, 68540, 
    68541, 68542, 68543, 68544, 68545, 68546, 68547, 68548, 68549, 68550, 
    68551, 68552, 68553, 68554, 68555, 68556, 68557, 68558, 68559, 68560, 
    68561, 68562, 68563, 68564, 68565, 68566, 68567, 68568, 68569, 68570, 
    68571, 68572, 68573, 68574, 68575, 68576, 68577, 68578, 68579, 68580, 
    68581, 68582, 68583, 68584, 68585, 68586, 68587, 68588, 68589, 68590, 
    68591, 68592, 68593, 68594, 68595, 68596, 68597, 68598, 68599, 68600, 
    68601, 68602, 68603, 68604, 68605, 68606, 68607, 68608, 68609, 68610, 
    68611, 68612, 68613, 68614, 68615, 68616, 68617, 68618, 68619, 68620, 
    68621, 68622, 68623, 68624, 68625, 68626, 68627, 68628, 68629, 68630, 
    68631, 68632, 68633, 68634, 68635, 68636, 68637, 68638, 68639, 68640, 
    68641, 68642, 68643, 68644, 68645, 68646, 68647, 68648, 68649, 68650, 
    68651, 68652, 68653, 68654, 68655, 68656, 68657, 68658, 68659, 68660, 
    68661, 68662, 68663, 68664, 68665, 68666, 68667, 68668, 68669, 68670, 
    68671, 68672, 68673, 68674, 68675, 68676, 68677, 68678, 68679, 68680, 
    68681, 68682, 68683, 68684, 68685, 68686, 68687, 68688, 68689, 68690, 
    68691, 68692, 68693, 68694, 68695, 68696, 68697, 68698, 68699, 68700, 
    68701, 68702, 68703, 68704, 68705, 68706, 68707, 68708, 68709, 68710, 
    68711, 68712, 68713, 68714, 68715, 68716, 68717, 68718, 68719, 68720, 
    68721, 68722, 68723, 68724, 68725, 68726, 68727, 68728, 68729, 68730, 
    68731, 68732, 68733, 68734, 68735, 68736, 68737, 68738, 68739, 68740, 
    68741, 68742, 68743, 68744, 68745, 68746, 68747, 68748, 68749, 68750, 
    68751, 68752, 68753, 68754, 68755, 68756, 68757, 68758, 68759, 68760, 
    68761, 68762, 68763, 68764, 68765, 68766, 68767, 68768, 68769, 68770, 
    68771, 68772, 68773, 68774, 68775, 68776, 68777, 68778, 68779, 68780, 
    68781, 68782, 68783, 68784, 68785, 68786, 68787, 68788, 68789, 68790, 
    68791, 68792, 68793, 68794, 68795, 68796, 68797, 68798, 68799, 68800, 
    68801, 68802, 68803, 68804, 68805, 68806, 68807, 68808, 68809, 68810, 
    68811, 68812, 68813, 68814, 68815, 68816, 68817, 68818, 68819, 68820, 
    68821, 68822, 68823, 68824, 68825, 68826, 68827, 68828, 68829, 68830, 
    68831, 68832, 68833, 68834, 68835, 68836, 68837, 68838, 68839, 68840, 
    68841, 68842, 68843, 68844, 68845, 68846, 68847, 68848, 68849, 68850, 
    68851, 68852, 68853, 68854, 68855, 68856, 68857, 68858, 68859, 68860, 
    68861, 68862, 68863, 68864, 68865, 68866, 68867, 68868, 68869, 68870, 
    68871, 68872, 68873, 68874, 68875, 68876, 68877, 68878, 68879, 68880, 
    68881, 68882, 68883, 68884, 68885, 68886, 68887, 68888, 68889, 68890, 
    68891, 68892, 68893, 68894, 68895, 68896, 68897, 68898, 68899, 68900, 
    68901, 68902, 68903, 68904, 68905, 68906, 68907, 68908, 68909, 68910, 
    68911, 68912, 68913, 68914, 68915, 68916, 68917, 68918, 68919, 68920, 
    68921, 68922, 68923, 68924, 68925, 68926, 68927, 68928, 68929, 68930, 
    68931, 68932, 68933, 68934, 68935, 68936, 68937, 68938, 68939, 68940, 
    68941, 68942, 68943, 68944, 68945, 68946, 68947, 68948, 68949, 68950, 
    68951, 68952, 68953, 68954, 68955, 68956, 68957, 68958, 68959, 68960, 
    68961, 68962, 68963, 68964, 68965, 68966, 68967, 68968, 68969, 68970, 
    68971, 68972, 68973, 68974, 68975, 68976, 68977, 68978, 68979, 68980, 
    68981, 68982, 68983, 68984, 68985, 68986, 68987, 68988, 68989, 68990, 
    68991, 68992, 68993, 68994, 68995, 68996, 68997, 68998, 68999, 69000, 
    69001, 69002, 69003, 69004, 69005, 69006, 69007, 69008, 69009, 69010, 
    69011, 69012, 69013, 69014, 69015, 69016, 69017, 69018, 69019, 69020, 
    69021, 69022, 69023, 69024, 69025, 69026, 69027, 69028, 69029, 69030, 
    69031, 69032, 69033, 69034, 69035, 69036, 69037, 69038, 69039, 69040, 
    69041, 69042, 69043, 69044, 69045, 69046, 69047, 69048, 69049, 69050, 
    69051, 69052, 69053, 69054, 69055, 69056, 69057, 69058, 69059, 69060, 
    69061, 69062, 69063, 69064, 69065, 69066, 69067, 69068, 69069, 69070, 
    69071, 69072, 69073, 69074, 69075, 69076, 69077, 69078, 69079, 69080, 
    69081, 69082, 69083, 69084, 69085, 69086, 69087, 69088, 69089, 69090, 
    69091, 69092, 69093, 69094, 69095, 69096, 69097, 69098, 69099, 69100, 
    69101, 69102, 69103, 69104, 69105, 69106, 69107, 69108, 69109, 69110, 
    69111, 69112, 69113, 69114, 69115, 69116, 69117, 69118, 69119, 69120, 
    69121, 69122, 69123, 69124, 69125, 69126, 69127, 69128, 69129, 69130, 
    69131, 69132, 69133, 69134, 69135, 69136, 69137, 69138, 69139, 69140, 
    69141, 69142, 69143, 69144, 69145, 69146, 69147, 69148, 69149, 69150, 
    69151, 69152, 69153, 69154, 69155, 69156, 69157, 69158, 69159, 69160, 
    69161, 69162, 69163, 69164, 69165, 69166, 69167, 69168, 69169, 69170, 
    69171, 69172, 69173, 69174, 69175, 69176, 69177, 69178, 69179, 69180, 
    69181, 69182, 69183, 69184, 69185, 69186, 69187, 69188, 69189, 69190, 
    69191, 69192, 69193, 69194, 69195, 69196, 69197, 69198, 69199, 69200, 
    69201, 69202, 69203, 69204, 69205, 69206, 69207, 69208, 69209, 69210, 
    69211, 69212, 69213, 69214, 69215, 69216, 69217, 69218, 69219, 69220, 
    69221, 69222, 69223, 69224, 69225, 69226, 69227, 69228, 69229, 69230, 
    69231, 69232, 69233, 69234, 69235, 69236, 69237, 69238, 69239, 69240, 
    69241, 69242, 69243, 69244, 69245, 69246, 69247, 69248, 69249, 69250, 
    69251, 69252, 69253, 69254, 69255, 69256, 69257, 69258, 69259, 69260, 
    69261, 69262, 69263, 69264, 69265, 69266, 69267, 69268, 69269, 69270, 
    69271, 69272, 69273, 69274, 69275, 69276, 69277, 69278, 69279, 69280, 
    69281, 69282, 69283, 69284, 69285, 69286, 69287, 69288, 69289, 69290, 
    69291, 69292, 69293, 69294, 69295, 69296, 69297, 69298, 69299, 69300, 
    69301, 69302, 69303, 69304, 69305, 69306, 69307, 69308, 69309, 69310, 
    69311, 69312, 69313, 69314, 69315, 69316, 69317, 69318, 69319, 69320, 
    69321, 69322, 69323, 69324, 69325, 69326, 69327, 69328, 69329, 69330, 
    69331, 69332, 69333, 69334, 69335, 69336, 69337, 69338, 69339, 69340, 
    69341, 69342, 69343, 69344, 69345, 69346, 69347, 69348, 69349, 69350, 
    69351, 69352, 69353, 69354, 69355, 69356, 69357, 69358, 69359, 69360, 
    69361, 69362, 69363, 69364, 69365, 69366, 69367, 69368, 69369, 69370, 
    69371, 69372, 69373, 69374, 69375, 69376, 69377, 69378, 69379, 69380, 
    69381, 69382, 69383, 69384, 69385, 69386, 69387, 69388, 69389, 69390, 
    69391, 69392, 69393, 69394, 69395, 69396, 69397, 69398, 69399, 69400, 
    69401, 69402, 69403, 69404, 69405, 69406, 69407, 69408, 69409, 69410, 
    69411, 69412, 69413, 69414, 69415, 69416, 69417, 69418, 69419, 69420, 
    69421, 69422, 69423, 69424, 69425, 69426, 69427, 69428, 69429, 69430, 
    69431, 69432, 69433, 69434, 69435, 69436, 69437, 69438, 69439, 69440, 
    69441, 69442, 69443, 69444, 69445, 69446, 69447, 69448, 69449, 69450, 
    69451, 69452, 69453, 69454, 69455, 69456, 69457, 69458, 69459, 69460, 
    69461, 69462, 69463, 69464, 69465, 69466, 69467, 69468, 69469, 69470, 
    69471, 69472, 69473, 69474, 69475, 69476, 69477, 69478, 69479, 69480, 
    69481, 69482, 69483, 69484, 69485, 69486, 69487, 69488, 69489, 69490, 
    69491, 69492, 69493, 69494, 69495, 69496, 69497, 69498, 69499, 69500, 
    69501, 69502, 69503, 69504, 69505, 69506, 69507, 69508, 69509, 69510, 
    69511, 69512, 69513, 69514, 69515, 69516, 69517, 69518, 69519, 69520, 
    69521, 69522, 69523, 69524, 69525, 69526, 69527, 69528, 69529, 69530, 
    69531, 69532, 69533, 69534, 69535, 69536, 69537, 69538, 69539, 69540, 
    69541, 69542, 69543, 69544, 69545, 69546, 69547, 69548, 69549, 69550, 
    69551, 69552, 69553, 69554, 69555, 69556, 69557, 69558, 69559, 69560, 
    69561, 69562, 69563, 69564, 69565, 69566, 69567, 69568, 69569, 69570, 
    69571, 69572, 69573, 69574, 69575, 69576, 69577, 69578, 69579, 69580, 
    69581, 69582, 69583, 69584, 69585, 69586, 69587, 69588, 69589, 69590, 
    69591, 69592, 69593, 69594, 69595, 69596, 69597, 69598, 69599, 69600, 
    69601, 69602, 69603, 69604, 69605, 69606, 69607, 69608, 69609, 69610, 
    69611, 69612, 69613, 69614, 69615, 69616, 69617, 69618, 69619, 69620, 
    69621, 69622, 69623, 69624, 69625, 69626, 69627, 69628, 69629, 69630, 
    69631, 69632, 69633, 69634, 69635, 69636, 69637, 69638, 69639, 69640, 
    69641, 69642, 69643, 69644, 69645, 69646, 69647, 69648, 69649, 69650, 
    69651, 69652, 69653, 69654, 69655, 69656, 69657, 69658, 69659, 69660, 
    69661, 69662, 69663, 69664, 69665, 69666, 69667, 69668, 69669, 69670, 
    69671, 69672, 69673, 69674, 69675, 69676, 69677, 69678, 69679, 69680, 
    69681, 69682, 69683, 69684, 69685, 69686, 69687, 69688, 69689, 69690, 
    69691, 69692, 69693, 69694, 69695, 69696, 69697, 69698, 69699, 69700, 
    69701, 69702, 69703, 69704, 69705, 69706, 69707, 69708, 69709, 69710, 
    69711, 69712, 69713, 69714, 69715, 69716, 69717, 69718, 69719, 69720, 
    69721, 69722, 69723, 69724, 69725, 69726, 69727, 69728, 69729, 69730, 
    69731, 69732, 69733, 69734, 69735, 69736, 69737, 69738, 69739, 69740, 
    69741, 69742, 69743, 69744, 69745, 69746, 69747, 69748, 69749, 69750, 
    69751, 69752, 69753, 69754, 69755, 69756, 69757, 69758, 69759, 69760, 
    69761, 69762, 69763, 69764, 69765, 69766, 69767, 69768, 69769, 69770, 
    69771, 69772, 69773, 69774, 69775, 69776, 69777, 69778, 69779, 69780, 
    69781, 69782, 69783, 69784, 69785, 69786, 69787, 69788, 69789, 69790, 
    69791, 69792, 69793, 69794, 69795, 69796, 69797, 69798, 69799, 69800, 
    69801, 69802, 69803, 69804, 69805, 69806, 69807, 69808, 69809, 69810, 
    69811, 69812, 69813, 69814, 69815, 69816, 69817, 69818, 69819, 69820, 
    69821, 69822, 69823, 69824, 69825, 69826, 69827, 69828, 69829, 69830, 
    69831, 69832, 69833, 69834, 69835, 69836, 69837, 69838, 69839, 69840, 
    69841, 69842, 69843, 69844, 69845, 69846, 69847, 69848, 69849, 69850, 
    69851, 69852, 69853, 69854, 69855, 69856, 69857, 69858, 69859, 69860, 
    69861, 69862, 69863, 69864, 69865, 69866, 69867, 69868, 69869, 69870, 
    69871, 69872, 69873, 69874, 69875, 69876, 69877, 69878, 69879, 69880, 
    69881, 69882, 69883, 69884, 69885, 69886, 69887, 69888, 69889, 69890, 
    69891, 69892, 69893, 69894, 69895, 69896, 69897, 69898, 69899, 69900, 
    69901, 69902, 69903, 69904, 69905, 69906, 69907, 69908, 69909, 69910, 
    69911, 69912, 69913, 69914, 69915, 69916, 69917, 69918, 69919, 69920, 
    69921, 69922, 69923, 69924, 69925, 69926, 69927, 69928, 69929, 69930, 
    69931, 69932, 69933, 69934, 69935, 69936, 69937, 69938, 69939, 69940, 
    69941, 69942, 69943, 69944, 69945, 69946, 69947, 69948, 69949, 69950, 
    69951, 69952, 69953, 69954, 69955, 69956, 69957, 69958, 69959, 69960, 
    69961, 69962, 69963, 69964, 69965, 69966, 69967, 69968, 69969, 69970, 
    69971, 69972, 69973, 69974, 69975, 69976, 69977, 69978, 69979, 69980, 
    69981, 69982, 69983, 69984, 69985, 69986, 69987, 69988, 69989, 69990, 
    69991, 69992, 69993, 69994, 69995, 69996, 69997, 69998, 69999, 70000, 
    70001, 70002, 70003, 70004, 70005, 70006, 70007, 70008, 70009, 70010, 
    70011, 70012, 70013, 70014, 70015, 70016, 70017, 70018, 70019, 70020, 
    70021, 70022, 70023, 70024, 70025, 70026, 70027, 70028, 70029, 70030, 
    70031, 70032, 70033, 70034, 70035, 70036, 70037, 70038, 70039, 70040, 
    70041, 70042, 70043, 70044, 70045, 70046, 70047, 70048, 70049, 70050, 
    70051, 70052, 70053, 70054, 70055, 70056, 70057, 70058, 70059, 70060, 
    70061, 70062, 70063, 70064, 70065, 70066, 70067, 70068, 70069, 70070, 
    70071, 70072, 70073, 70074, 70075, 70076, 70077, 70078, 70079, 70080, 
    70081, 70082, 70083, 70084, 70085, 70086, 70087, 70088, 70089, 70090, 
    70091, 70092, 70093, 70094, 70095, 70096, 70097, 70098, 70099, 70100, 
    70101, 70102, 70103, 70104, 70105, 70106, 70107, 70108, 70109, 70110, 
    70111, 70112, 70113, 70114, 70115, 70116, 70117, 70118, 70119, 70120, 
    70121, 70122, 70123, 70124, 70125, 70126, 70127, 70128, 70129, 70130, 
    70131, 70132, 70133, 70134, 70135, 70136, 70137, 70138, 70139, 70140, 
    70141, 70142, 70143, 70144, 70145, 70146, 70147, 70148, 70149, 70150, 
    70151, 70152, 70153, 70154, 70155, 70156, 70157, 70158, 70159, 70160, 
    70161, 70162, 70163, 70164, 70165, 70166, 70167, 70168, 70169, 70170, 
    70171, 70172, 70173, 70174, 70175, 70176, 70177, 70178, 70179, 70180, 
    70181, 70182, 70183, 70184, 70185, 70186, 70187, 70188, 70189, 70190, 
    70191, 70192, 70193, 70194, 70195, 70196, 70197, 70198, 70199, 70200, 
    70201, 70202, 70203, 70204, 70205, 70206, 70207, 70208, 70209, 70210, 
    70211, 70212, 70213, 70214, 70215, 70216, 70217, 70218, 70219, 70220, 
    70221, 70222, 70223, 70224, 70225, 70226, 70227, 70228, 70229, 70230, 
    70231, 70232, 70233, 70234, 70235, 70236, 70237, 70238, 70239, 70240, 
    70241, 70242, 70243, 70244, 70245, 70246, 70247, 70248, 70249, 70250, 
    70251, 70252, 70253, 70254, 70255, 70256, 70257, 70258, 70259, 70260, 
    70261, 70262, 70263, 70264, 70265, 70266, 70267, 70268, 70269, 70270, 
    70271, 70272, 70273, 70274, 70275, 70276, 70277, 70278, 70279, 70280, 
    70281, 70282, 70283, 70284, 70285, 70286, 70287, 70288, 70289, 70290, 
    70291, 70292, 70293, 70294, 70295, 70296, 70297, 70298, 70299, 70300, 
    70301, 70302, 70303, 70304, 70305, 70306, 70307, 70308, 70309, 70310, 
    70311, 70312, 70313, 70314, 70315, 70316, 70317, 70318, 70319, 70320, 
    70321, 70322, 70323, 70324, 70325, 70326, 70327, 70328, 70329, 70330, 
    70331, 70332, 70333, 70334, 70335, 70336, 70337, 70338, 70339, 70340, 
    70341, 70342, 70343, 70344, 70345, 70346, 70347, 70348, 70349, 70350, 
    70351, 70352, 70353, 70354, 70355, 70356, 70357, 70358, 70359, 70360, 
    70361, 70362, 70363, 70364, 70365, 70366, 70367, 70368, 70369, 70370, 
    70371, 70372, 70373, 70374, 70375, 70376, 70377, 70378, 70379, 70380, 
    70381, 70382, 70383, 70384, 70385, 70386, 70387, 70388, 70389, 70390, 
    70391, 70392, 70393, 70394, 70395, 70396, 70397, 70398, 70399, 70400, 
    70401, 70402, 70403, 70404, 70405, 70406, 70407, 70408, 70409, 70410, 
    70411, 70412, 70413, 70414, 70415, 70416, 70417, 70418, 70419, 70420, 
    70421, 70422, 70423, 70424, 70425, 70426, 70427, 70428, 70429, 70430, 
    70431, 70432, 70433, 70434, 70435, 70436, 70437, 70438, 70439, 70440, 
    70441, 70442, 70443, 70444, 70445, 70446, 70447, 70448, 70449, 70450, 
    70451, 70452, 70453, 70454, 70455, 70456, 70457, 70458, 70459, 70460, 
    70461, 70462, 70463, 70464, 70465, 70466, 70467, 70468, 70469, 70470, 
    70471, 70472, 70473, 70474, 70475, 70476, 70477, 70478, 70479, 70480, 
    70481, 70482, 70483, 70484, 70485, 70486, 70487, 70488, 70489, 70490, 
    70491, 70492, 70493, 70494, 70495, 70496, 70497, 70498, 70499, 70500, 
    70501, 70502, 70503, 70504, 70505, 70506, 70507, 70508, 70509, 70510, 
    70511, 70512, 70513, 70514, 70515, 70516, 70517, 70518, 70519, 70520, 
    70521, 70522, 70523, 70524, 70525, 70526, 70527, 70528, 70529, 70530, 
    70531, 70532, 70533, 70534, 70535, 70536, 70537, 70538, 70539, 70540, 
    70541, 70542, 70543, 70544, 70545, 70546, 70547, 70548, 70549, 70550, 
    70551, 70552, 70553, 70554, 70555, 70556, 70557, 70558, 70559, 70560, 
    70561, 70562, 70563, 70564, 70565, 70566, 70567, 70568, 70569, 70570, 
    70571, 70572, 70573, 70574, 70575, 70576, 70577, 70578, 70579, 70580, 
    70581, 70582, 70583, 70584, 70585, 70586, 70587, 70588, 70589, 70590, 
    70591, 70592, 70593, 70594, 70595, 70596, 70597, 70598, 70599, 70600, 
    70601, 70602, 70603, 70604, 70605, 70606, 70607, 70608, 70609, 70610, 
    70611, 70612, 70613, 70614, 70615, 70616, 70617, 70618, 70619, 70620, 
    70621, 70622, 70623, 70624, 70625, 70626, 70627, 70628, 70629, 70630, 
    70631, 70632, 70633, 70634, 70635, 70636, 70637, 70638, 70639, 70640, 
    70641, 70642, 70643, 70644, 70645, 70646, 70647, 70648, 70649, 70650, 
    70651, 70652, 70653, 70654, 70655, 70656, 70657, 70658, 70659, 70660, 
    70661, 70662, 70663, 70664, 70665, 70666, 70667, 70668, 70669, 70670, 
    70671, 70672, 70673, 70674, 70675, 70676, 70677, 70678, 70679, 70680, 
    70681, 70682, 70683, 70684, 70685, 70686, 70687, 70688, 70689, 70690, 
    70691, 70692, 70693, 70694, 70695, 70696, 70697, 70698, 70699, 70700, 
    70701, 70702, 70703, 70704, 70705, 70706, 70707, 70708, 70709, 70710, 
    70711, 70712, 70713, 70714, 70715, 70716, 70717, 70718, 70719, 70720, 
    70721, 70722, 70723, 70724, 70725, 70726, 70727, 70728, 70729, 70730, 
    70731, 70732, 70733, 70734, 70735, 70736, 70737, 70738, 70739, 70740, 
    70741, 70742, 70743, 70744, 70745, 70746, 70747, 70748, 70749, 70750, 
    70751, 70752, 70753, 70754, 70755, 70756, 70757, 70758, 70759, 70760, 
    70761, 70762, 70763, 70764, 70765, 70766, 70767, 70768, 70769, 70770, 
    70771, 70772, 70773, 70774, 70775, 70776, 70777, 70778, 70779, 70780, 
    70781, 70782, 70783, 70784, 70785, 70786, 70787, 70788, 70789, 70790, 
    70791, 70792, 70793, 70794, 70795, 70796, 70797, 70798, 70799, 70800, 
    70801, 70802, 70803, 70804, 70805, 70806, 70807, 70808, 70809, 70810, 
    70811, 70812, 70813, 70814, 70815, 70816, 70817, 70818, 70819, 70820, 
    70821, 70822, 70823, 70824, 70825, 70826, 70827, 70828, 70829, 70830, 
    70831, 70832, 70833, 70834, 70835, 70836, 70837, 70838, 70839, 70840, 
    70841, 70842, 70843, 70844, 70845, 70846, 70847, 70848, 70849, 70850, 
    70851, 70852, 70853, 70854, 70855, 70856, 70857, 70858, 70859, 70860, 
    70861, 70862, 70863, 70864, 70865, 70866, 70867, 70868, 70869, 70870, 
    70871, 70872, 70873, 70874, 70875, 70876, 70877, 70878, 70879, 70880, 
    70881, 70882, 70883, 70884, 70885, 70886, 70887, 70888, 70889, 70890, 
    70891, 70892, 70893, 70894, 70895, 70896, 70897, 70898, 70899, 70900, 
    70901, 70902, 70903, 70904, 70905, 70906, 70907, 70908, 70909, 70910, 
    70911, 70912, 70913, 70914, 70915, 70916, 70917, 70918, 70919, 70920, 
    70921, 70922, 70923, 70924, 70925, 70926, 70927, 70928, 70929, 70930, 
    70931, 70932, 70933, 70934, 70935, 70936, 70937, 70938, 70939, 70940, 
    70941, 70942, 70943, 70944, 70945, 70946, 70947, 70948, 70949, 70950, 
    70951, 70952, 70953, 70954, 70955, 70956, 70957, 70958, 70959, 70960, 
    70961, 70962, 70963, 70964, 70965, 70966, 70967, 70968, 70969, 70970, 
    70971, 70972, 70973, 70974, 70975, 70976, 70977, 70978, 70979, 70980, 
    70981, 70982, 70983, 70984, 70985, 70986, 70987, 70988, 70989, 70990, 
    70991, 70992, 70993, 70994, 70995, 70996, 70997, 70998, 70999, 71000, 
    71001, 71002, 71003, 71004, 71005, 71006, 71007, 71008, 71009, 71010, 
    71011, 71012, 71013, 71014, 71015, 71016, 71017, 71018, 71019, 71020, 
    71021, 71022, 71023, 71024, 71025, 71026, 71027, 71028, 71029, 71030, 
    71031, 71032, 71033, 71034, 71035, 71036, 71037, 71038, 71039, 71040, 
    71041, 71042, 71043, 71044, 71045, 71046, 71047, 71048, 71049, 71050, 
    71051, 71052, 71053, 71054, 71055, 71056, 71057, 71058, 71059, 71060, 
    71061, 71062, 71063, 71064, 71065, 71066, 71067, 71068, 71069, 71070, 
    71071, 71072, 71073, 71074, 71075, 71076, 71077, 71078, 71079, 71080, 
    71081, 71082, 71083, 71084, 71085, 71086, 71087, 71088, 71089, 71090, 
    71091, 71092, 71093, 71094, 71095, 71096, 71097, 71098, 71099, 71100, 
    71101, 71102, 71103, 71104, 71105, 71106, 71107, 71108, 71109, 71110, 
    71111, 71112, 71113, 71114, 71115, 71116, 71117, 71118, 71119, 71120, 
    71121, 71122, 71123, 71124, 71125, 71126, 71127, 71128, 71129, 71130, 
    71131, 71132, 71133, 71134, 71135, 71136, 71137, 71138, 71139, 71140, 
    71141, 71142, 71143, 71144, 71145, 71146, 71147, 71148, 71149, 71150, 
    71151, 71152, 71153, 71154, 71155, 71156, 71157, 71158, 71159, 71160, 
    71161, 71162, 71163, 71164, 71165, 71166, 71167, 71168, 71169, 71170, 
    71171, 71172, 71173, 71174, 71175, 71176, 71177, 71178, 71179, 71180, 
    71181, 71182, 71183, 71184, 71185, 71186, 71187, 71188, 71189, 71190, 
    71191, 71192, 71193, 71194, 71195, 71196, 71197, 71198, 71199, 71200, 
    71201, 71202, 71203, 71204, 71205, 71206, 71207, 71208, 71209, 71210, 
    71211, 71212, 71213, 71214, 71215, 71216, 71217, 71218, 71219, 71220, 
    71221, 71222, 71223, 71224, 71225, 71226, 71227, 71228, 71229, 71230, 
    71231, 71232, 71233, 71234, 71235, 71236, 71237, 71238, 71239, 71240, 
    71241, 71242, 71243, 71244, 71245, 71246, 71247, 71248, 71249, 71250, 
    71251, 71252, 71253, 71254, 71255, 71256, 71257, 71258, 71259, 71260, 
    71261, 71262, 71263, 71264, 71265, 71266, 71267, 71268, 71269, 71270, 
    71271, 71272, 71273, 71274, 71275, 71276, 71277, 71278, 71279, 71280, 
    71281, 71282, 71283, 71284, 71285, 71286, 71287, 71288, 71289, 71290, 
    71291, 71292, 71293, 71294, 71295, 71296, 71297, 71298, 71299, 71300, 
    71301, 71302, 71303, 71304, 71305, 71306, 71307, 71308, 71309, 71310, 
    71311, 71312, 71313, 71314, 71315, 71316, 71317, 71318, 71319, 71320, 
    71321, 71322, 71323, 71324, 71325, 71326, 71327, 71328, 71329, 71330, 
    71331, 71332, 71333, 71334, 71335, 71336, 71337, 71338, 71339, 71340, 
    71341, 71342, 71343, 71344, 71345, 71346, 71347, 71348, 71349, 71350, 
    71351, 71352, 71353, 71354, 71355, 71356, 71357, 71358, 71359, 71360, 
    71361, 71362, 71363, 71364, 71365, 71366, 71367, 71368, 71369, 71370, 
    71371, 71372, 71373, 71374, 71375, 71376, 71377, 71378, 71379, 71380, 
    71381, 71382, 71383, 71384, 71385, 71386, 71387, 71388, 71389, 71390, 
    71391, 71392, 71393, 71394, 71395, 71396, 71397, 71398, 71399, 71400, 
    71401, 71402, 71403, 71404, 71405, 71406, 71407, 71408, 71409, 71410, 
    71411, 71412, 71413, 71414, 71415, 71416, 71417, 71418, 71419, 71420, 
    71421, 71422, 71423, 71424, 71425, 71426, 71427, 71428, 71429, 71430, 
    71431, 71432, 71433, 71434, 71435, 71436, 71437, 71438, 71439, 71440, 
    71441, 71442, 71443, 71444, 71445, 71446, 71447, 71448, 71449, 71450, 
    71451, 71452, 71453, 71454, 71455, 71456, 71457, 71458, 71459, 71460, 
    71461, 71462, 71463, 71464, 71465, 71466, 71467, 71468, 71469, 71470, 
    71471, 71472, 71473, 71474, 71475, 71476, 71477, 71478, 71479, 71480, 
    71481, 71482, 71483, 71484, 71485, 71486, 71487, 71488, 71489, 71490, 
    71491, 71492, 71493, 71494, 71495, 71496, 71497, 71498, 71499, 71500, 
    71501, 71502, 71503, 71504, 71505, 71506, 71507, 71508, 71509, 71510, 
    71511, 71512, 71513, 71514, 71515, 71516, 71517, 71518, 71519, 71520, 
    71521, 71522, 71523, 71524, 71525, 71526, 71527, 71528, 71529, 71530, 
    71531, 71532, 71533, 71534, 71535, 71536, 71537, 71538, 71539, 71540, 
    71541, 71542, 71543, 71544, 71545, 71546, 71547, 71548, 71549, 71550, 
    71551, 71552, 71553, 71554, 71555, 71556, 71557, 71558, 71559, 71560, 
    71561, 71562, 71563, 71564, 71565, 71566, 71567, 71568, 71569, 71570, 
    71571, 71572, 71573, 71574, 71575, 71576, 71577, 71578, 71579, 71580, 
    71581, 71582, 71583, 71584, 71585, 71586, 71587, 71588, 71589, 71590, 
    71591, 71592, 71593, 71594, 71595, 71596, 71597, 71598, 71599, 71600, 
    71601, 71602, 71603, 71604, 71605, 71606, 71607, 71608, 71609, 71610, 
    71611, 71612, 71613, 71614, 71615, 71616, 71617, 71618, 71619, 71620, 
    71621, 71622, 71623, 71624, 71625, 71626, 71627, 71628, 71629, 71630, 
    71631, 71632, 71633, 71634, 71635, 71636, 71637, 71638, 71639, 71640, 
    71641, 71642, 71643, 71644, 71645, 71646, 71647, 71648, 71649, 71650, 
    71651, 71652, 71653, 71654, 71655, 71656, 71657, 71658, 71659, 71660, 
    71661, 71662, 71663, 71664, 71665, 71666, 71667, 71668, 71669, 71670, 
    71671, 71672, 71673, 71674, 71675, 71676, 71677, 71678, 71679, 71680, 
    71681, 71682, 71683, 71684, 71685, 71686, 71687, 71688, 71689, 71690, 
    71691, 71692, 71693, 71694, 71695, 71696, 71697, 71698, 71699, 71700, 
    71701, 71702, 71703, 71704, 71705, 71706, 71707, 71708, 71709, 71710, 
    71711, 71712, 71713, 71714, 71715, 71716, 71717, 71718, 71719, 71720, 
    71721, 71722, 71723, 71724, 71725, 71726, 71727, 71728, 71729, 71730, 
    71731, 71732, 71733, 71734, 71735, 71736, 71737, 71738, 71739, 71740, 
    71741, 71742, 71743, 71744, 71745, 71746, 71747, 71748, 71749, 71750, 
    71751, 71752, 71753, 71754, 71755, 71756, 71757, 71758, 71759, 71760, 
    71761, 71762, 71763, 71764, 71765, 71766, 71767, 71768, 71769, 71770, 
    71771, 71772, 71773, 71774, 71775, 71776, 71777, 71778, 71779, 71780, 
    71781, 71782, 71783, 71784, 71785, 71786, 71787, 71788, 71789, 71790, 
    71791, 71792, 71793, 71794, 71795, 71796, 71797, 71798, 71799, 71800, 
    71801, 71802, 71803, 71804, 71805, 71806, 71807, 71808, 71809, 71810, 
    71811, 71812, 71813, 71814, 71815, 71816, 71817, 71818, 71819, 71820, 
    71821, 71822, 71823, 71824, 71825, 71826, 71827, 71828, 71829, 71830, 
    71831, 71832, 71833, 71834, 71835, 71836, 71837, 71838, 71839, 71840, 
    71841, 71842, 71843, 71844, 71845, 71846, 71847, 71848, 71849, 71850, 
    71851, 71852, 71853, 71854, 71855, 71856, 71857, 71858, 71859, 71860, 
    71861, 71862, 71863, 71864, 71865, 71866, 71867, 71868, 71869, 71870, 
    71871, 71872, 71873, 71874, 71875, 71876, 71877, 71878, 71879, 71880, 
    71881, 71882, 71883, 71884, 71885, 71886, 71887, 71888, 71889, 71890, 
    71891, 71892, 71893, 71894, 71895, 71896, 71897, 71898, 71899, 71900, 
    71901, 71902, 71903, 71904, 71905, 71906, 71907, 71908, 71909, 71910, 
    71911, 71912, 71913, 71914, 71915, 71916, 71917, 71918, 71919, 71920, 
    71921, 71922, 71923, 71924, 71925, 71926, 71927, 71928, 71929, 71930, 
    71931, 71932, 71933, 71934, 71935, 71936, 71937, 71938, 71939, 71940, 
    71941, 71942, 71943, 71944, 71945, 71946, 71947, 71948, 71949, 71950, 
    71951, 71952, 71953, 71954, 71955, 71956, 71957, 71958, 71959, 71960, 
    71961, 71962, 71963, 71964, 71965, 71966, 71967, 71968, 71969, 71970, 
    71971, 71972, 71973, 71974, 71975, 71976, 71977, 71978, 71979, 71980, 
    71981, 71982, 71983, 71984, 71985, 71986, 71987, 71988, 71989, 71990, 
    71991, 71992, 71993, 71994, 71995, 71996, 71997, 71998, 71999, 72000, 
    72001, 72002, 72003, 72004, 72005, 72006, 72007, 72008, 72009, 72010, 
    72011, 72012, 72013, 72014, 72015, 72016, 72017, 72018, 72019, 72020, 
    72021, 72022, 72023, 72024, 72025, 72026, 72027, 72028, 72029, 72030, 
    72031, 72032, 72033, 72034, 72035, 72036, 72037, 72038, 72039, 72040, 
    72041, 72042, 72043, 72044, 72045, 72046, 72047, 72048, 72049, 72050, 
    72051, 72052, 72053, 72054, 72055, 72056, 72057, 72058, 72059, 72060, 
    72061, 72062, 72063, 72064, 72065, 72066, 72067, 72068, 72069, 72070, 
    72071, 72072, 72073, 72074, 72075, 72076, 72077, 72078, 72079, 72080, 
    72081, 72082, 72083, 72084, 72085, 72086, 72087, 72088, 72089, 72090, 
    72091, 72092, 72093, 72094, 72095, 72096, 72097, 72098, 72099, 72100, 
    72101, 72102, 72103, 72104, 72105, 72106, 72107, 72108, 72109, 72110, 
    72111, 72112, 72113, 72114, 72115, 72116, 72117, 72118, 72119, 72120, 
    72121, 72122, 72123, 72124, 72125, 72126, 72127, 72128, 72129, 72130, 
    72131, 72132, 72133, 72134, 72135, 72136, 72137, 72138, 72139, 72140, 
    72141, 72142, 72143, 72144, 72145, 72146, 72147, 72148, 72149, 72150, 
    72151, 72152, 72153, 72154, 72155, 72156, 72157, 72158, 72159, 72160, 
    72161, 72162, 72163, 72164, 72165, 72166, 72167, 72168, 72169, 72170, 
    72171, 72172, 72173, 72174, 72175, 72176, 72177, 72178, 72179, 72180, 
    72181, 72182, 72183, 72184, 72185, 72186, 72187, 72188, 72189, 72190, 
    72191, 72192, 72193, 72194, 72195, 72196, 72197, 72198, 72199, 72200, 
    72201, 72202, 72203, 72204, 72205, 72206, 72207, 72208, 72209, 72210, 
    72211, 72212, 72213, 72214, 72215, 72216, 72217, 72218, 72219, 72220, 
    72221, 72222, 72223, 72224, 72225, 72226, 72227, 72228, 72229, 72230, 
    72231, 72232, 72233, 72234, 72235, 72236, 72237, 72238, 72239, 72240, 
    72241, 72242, 72243, 72244, 72245, 72246, 72247, 72248, 72249, 72250, 
    72251, 72252, 72253, 72254, 72255, 72256, 72257, 72258, 72259, 72260, 
    72261, 72262, 72263, 72264, 72265, 72266, 72267, 72268, 72269, 72270, 
    72271, 72272, 72273, 72274, 72275, 72276, 72277, 72278, 72279, 72280, 
    72281, 72282, 72283, 72284, 72285, 72286, 72287, 72288, 72289, 72290, 
    72291, 72292, 72293, 72294, 72295, 72296, 72297, 72298, 72299, 72300, 
    72301, 72302, 72303, 72304, 72305, 72306, 72307, 72308, 72309, 72310, 
    72311, 72312, 72313, 72314, 72315, 72316, 72317, 72318, 72319, 72320, 
    72321, 72322, 72323, 72324, 72325, 72326, 72327, 72328, 72329, 72330, 
    72331, 72332, 72333, 72334, 72335, 72336, 72337, 72338, 72339, 72340, 
    72341, 72342, 72343, 72344, 72345, 72346, 72347, 72348, 72349, 72350, 
    72351, 72352, 72353, 72354, 72355, 72356, 72357, 72358, 72359, 72360, 
    72361, 72362, 72363, 72364, 72365, 72366, 72367, 72368, 72369, 72370, 
    72371, 72372, 72373, 72374, 72375, 72376, 72377, 72378, 72379, 72380, 
    72381, 72382, 72383, 72384, 72385, 72386, 72387, 72388, 72389, 72390, 
    72391, 72392, 72393, 72394, 72395, 72396, 72397, 72398, 72399, 72400, 
    72401, 72402, 72403, 72404, 72405, 72406, 72407, 72408, 72409, 72410, 
    72411, 72412, 72413, 72414, 72415, 72416, 72417, 72418, 72419, 72420, 
    72421, 72422, 72423, 72424, 72425, 72426, 72427, 72428, 72429, 72430, 
    72431, 72432, 72433, 72434, 72435, 72436, 72437, 72438, 72439, 72440, 
    72441, 72442, 72443, 72444, 72445, 72446, 72447, 72448, 72449, 72450, 
    72451, 72452, 72453, 72454, 72455, 72456, 72457, 72458, 72459, 72460, 
    72461, 72462, 72463, 72464, 72465, 72466, 72467, 72468, 72469, 72470, 
    72471, 72472, 72473, 72474, 72475, 72476, 72477, 72478, 72479, 72480, 
    72481, 72482, 72483, 72484, 72485, 72486, 72487, 72488, 72489, 72490, 
    72491, 72492, 72493, 72494, 72495, 72496, 72497, 72498, 72499, 72500, 
    72501, 72502, 72503, 72504, 72505, 72506, 72507, 72508, 72509, 72510, 
    72511, 72512, 72513, 72514, 72515, 72516, 72517, 72518, 72519, 72520, 
    72521, 72522, 72523, 72524, 72525, 72526, 72527, 72528, 72529, 72530, 
    72531, 72532, 72533, 72534, 72535, 72536, 72537, 72538, 72539, 72540, 
    72541, 72542, 72543, 72544, 72545, 72546, 72547, 72548, 72549, 72550, 
    72551, 72552, 72553, 72554, 72555, 72556, 72557, 72558, 72559, 72560, 
    72561, 72562, 72563, 72564, 72565, 72566, 72567, 72568, 72569, 72570, 
    72571, 72572, 72573, 72574, 72575, 72576, 72577, 72578, 72579, 72580, 
    72581, 72582, 72583, 72584, 72585, 72586, 72587, 72588, 72589, 72590, 
    72591, 72592, 72593, 72594, 72595, 72596, 72597, 72598, 72599, 72600, 
    72601, 72602, 72603, 72604, 72605, 72606, 72607, 72608, 72609, 72610, 
    72611, 72612, 72613, 72614, 72615, 72616, 72617, 72618, 72619, 72620, 
    72621, 72622, 72623, 72624, 72625, 72626, 72627, 72628, 72629, 72630, 
    72631, 72632, 72633, 72634, 72635, 72636, 72637, 72638, 72639, 72640, 
    72641, 72642, 72643, 72644, 72645, 72646, 72647, 72648, 72649, 72650, 
    72651, 72652, 72653, 72654, 72655, 72656, 72657, 72658, 72659, 72660, 
    72661, 72662, 72663, 72664, 72665, 72666, 72667, 72668, 72669, 72670, 
    72671, 72672, 72673, 72674, 72675, 72676, 72677, 72678, 72679, 72680, 
    72681, 72682, 72683, 72684, 72685, 72686, 72687, 72688, 72689, 72690, 
    72691, 72692, 72693, 72694, 72695, 72696, 72697, 72698, 72699, 72700, 
    72701, 72702, 72703, 72704, 72705, 72706, 72707, 72708, 72709, 72710, 
    72711, 72712, 72713, 72714, 72715, 72716, 72717, 72718, 72719, 72720, 
    72721, 72722, 72723, 72724, 72725, 72726, 72727, 72728, 72729, 72730, 
    72731, 72732, 72733, 72734, 72735, 72736, 72737, 72738, 72739, 72740, 
    72741, 72742, 72743, 72744, 72745, 72746, 72747, 72748, 72749, 72750, 
    72751, 72752, 72753, 72754, 72755, 72756, 72757, 72758, 72759, 72760, 
    72761, 72762, 72763, 72764, 72765, 72766, 72767, 72768, 72769, 72770, 
    72771, 72772, 72773, 72774, 72775, 72776, 72777, 72778, 72779, 72780, 
    72781, 72782, 72783, 72784, 72785, 72786, 72787, 72788, 72789, 72790, 
    72791, 72792, 72793, 72794, 72795, 72796, 72797, 72798, 72799, 72800, 
    72801, 72802, 72803, 72804, 72805, 72806, 72807, 72808, 72809, 72810, 
    72811, 72812, 72813, 72814, 72815, 72816, 72817, 72818, 72819, 72820, 
    72821, 72822, 72823, 72824, 72825, 72826, 72827, 72828, 72829, 72830, 
    72831, 72832, 72833, 72834, 72835, 72836, 72837, 72838, 72839, 72840, 
    72841, 72842, 72843, 72844, 72845, 72846, 72847, 72848, 72849, 72850, 
    72851, 72852, 72853, 72854, 72855, 72856, 72857, 72858, 72859, 72860, 
    72861, 72862, 72863, 72864, 72865, 72866, 72867, 72868, 72869, 72870, 
    72871, 72872, 72873, 72874, 72875, 72876, 72877, 72878, 72879, 72880, 
    72881, 72882, 72883, 72884, 72885, 72886, 72887, 72888, 72889, 72890, 
    72891, 72892, 72893, 72894, 72895, 72896, 72897, 72898, 72899, 72900, 
    72901, 72902, 72903, 72904, 72905, 72906, 72907, 72908, 72909, 72910, 
    72911, 72912, 72913, 72914, 72915, 72916, 72917, 72918, 72919, 72920, 
    72921, 72922, 72923, 72924, 72925, 72926, 72927, 72928, 72929, 72930, 
    72931, 72932, 72933, 72934, 72935, 72936, 72937, 72938, 72939, 72940, 
    72941, 72942, 72943, 72944, 72945, 72946, 72947, 72948, 72949, 72950, 
    72951, 72952, 72953, 72954, 72955, 72956, 72957, 72958, 72959, 72960, 
    72961, 72962, 72963, 72964, 72965, 72966, 72967, 72968, 72969, 72970, 
    72971, 72972, 72973, 72974, 72975, 72976, 72977, 72978, 72979, 72980, 
    72981, 72982, 72983, 72984, 72985, 72986, 72987, 72988, 72989, 72990, 
    72991, 72992, 72993, 72994, 72995, 72996, 72997, 72998, 72999, 73000, 
    73001, 73002, 73003, 73004, 73005, 73006, 73007, 73008, 73009, 73010, 
    73011, 73012, 73013, 73014, 73015, 73016, 73017, 73018, 73019, 73020, 
    73021, 73022, 73023, 73024, 73025, 73026, 73027, 73028, 73029, 73030, 
    73031, 73032, 73033, 73034, 73035, 73036, 73037, 73038, 73039, 73040, 
    73041, 73042, 73043, 73044, 73045, 73046, 73047, 73048, 73049, 73050, 
    73051, 73052, 73053, 73054, 73055, 73056, 73057, 73058, 73059, 73060, 
    73061, 73062, 73063, 73064, 73065, 73066, 73067, 73068, 73069, 73070, 
    73071, 73072, 73073, 73074, 73075, 73076, 73077, 73078, 73079, 73080, 
    73081, 73082, 73083, 73084, 73085, 73086, 73087, 73088, 73089, 73090, 
    73091, 73092, 73093, 73094, 73095, 73096, 73097, 73098, 73099, 73100, 
    73101, 73102, 73103, 73104, 73105, 73106, 73107, 73108, 73109, 73110, 
    73111, 73112, 73113, 73114, 73115, 73116, 73117, 73118, 73119, 73120, 
    73121, 73122, 73123, 73124, 73125, 73126, 73127, 73128, 73129, 73130, 
    73131, 73132, 73133, 73134, 73135, 73136, 73137, 73138, 73139, 73140, 
    73141, 73142, 73143, 73144, 73145, 73146, 73147, 73148, 73149, 73150, 
    73151, 73152, 73153, 73154, 73155, 73156, 73157, 73158, 73159, 73160, 
    73161, 73162, 73163, 73164, 73165, 73166, 73167, 73168, 73169, 73170, 
    73171, 73172, 73173, 73174, 73175, 73176, 73177, 73178, 73179, 73180, 
    73181, 73182, 73183, 73184, 73185, 73186, 73187, 73188, 73189, 73190, 
    73191, 73192, 73193, 73194, 73195, 73196, 73197, 73198, 73199, 73200, 
    73201, 73202, 73203, 73204, 73205, 73206, 73207, 73208, 73209, 73210, 
    73211, 73212, 73213, 73214, 73215, 73216, 73217, 73218, 73219, 73220, 
    73221, 73222, 73223, 73224, 73225, 73226, 73227, 73228, 73229, 73230, 
    73231, 73232, 73233, 73234, 73235, 73236, 73237, 73238, 73239, 73240, 
    73241, 73242, 73243, 73244, 73245, 73246, 73247, 73248, 73249, 73250, 
    73251, 73252, 73253, 73254, 73255, 73256, 73257, 73258, 73259, 73260, 
    73261, 73262, 73263, 73264, 73265, 73266, 73267, 73268, 73269, 73270, 
    73271, 73272, 73273, 73274, 73275, 73276, 73277, 73278, 73279, 73280, 
    73281, 73282, 73283, 73284, 73285, 73286, 73287, 73288, 73289, 73290, 
    73291, 73292, 73293, 73294, 73295, 73296, 73297, 73298, 73299, 73300, 
    73301, 73302, 73303, 73304, 73305, 73306, 73307, 73308, 73309, 73310, 
    73311, 73312, 73313, 73314, 73315, 73316, 73317, 73318, 73319, 73320, 
    73321, 73322, 73323, 73324, 73325, 73326, 73327, 73328, 73329, 73330, 
    73331, 73332, 73333, 73334, 73335, 73336, 73337, 73338, 73339, 73340, 
    73341, 73342, 73343, 73344, 73345, 73346, 73347, 73348, 73349, 73350, 
    73351, 73352, 73353, 73354, 73355, 73356, 73357, 73358, 73359, 73360, 
    73361, 73362, 73363, 73364, 73365, 73366, 73367, 73368, 73369, 73370, 
    73371, 73372, 73373, 73374, 73375, 73376, 73377, 73378, 73379, 73380, 
    73381, 73382, 73383, 73384, 73385, 73386, 73387, 73388, 73389, 73390, 
    73391, 73392, 73393, 73394, 73395, 73396, 73397, 73398, 73399, 73400, 
    73401, 73402, 73403, 73404, 73405, 73406, 73407, 73408, 73409, 73410, 
    73411, 73412, 73413, 73414, 73415, 73416, 73417, 73418, 73419, 73420, 
    73421, 73422, 73423, 73424, 73425, 73426, 73427, 73428, 73429, 73430, 
    73431, 73432, 73433, 73434, 73435, 73436, 73437, 73438, 73439, 73440, 
    73441, 73442, 73443, 73444, 73445, 73446, 73447, 73448, 73449, 73450, 
    73451, 73452, 73453, 73454, 73455, 73456, 73457, 73458, 73459, 73460, 
    73461, 73462, 73463, 73464, 73465, 73466, 73467, 73468, 73469, 73470, 
    73471, 73472, 73473, 73474, 73475, 73476, 73477, 73478, 73479, 73480, 
    73481, 73482, 73483, 73484, 73485, 73486, 73487, 73488, 73489, 73490, 
    73491, 73492, 73493, 73494, 73495, 73496, 73497, 73498, 73499, 73500, 
    73501, 73502, 73503, 73504, 73505, 73506, 73507, 73508, 73509, 73510, 
    73511, 73512, 73513, 73514, 73515, 73516, 73517, 73518, 73519, 73520, 
    73521, 73522, 73523, 73524, 73525, 73526, 73527, 73528, 73529, 73530, 
    73531, 73532, 73533, 73534, 73535, 73536, 73537, 73538, 73539, 73540, 
    73541, 73542, 73543, 73544, 73545, 73546, 73547, 73548, 73549, 73550, 
    73551, 73552, 73553, 73554, 73555, 73556, 73557, 73558, 73559, 73560, 
    73561, 73562, 73563, 73564, 73565, 73566, 73567, 73568, 73569, 73570, 
    73571, 73572, 73573, 73574, 73575, 73576, 73577, 73578, 73579, 73580, 
    73581, 73582, 73583, 73584, 73585, 73586, 73587, 73588, 73589, 73590, 
    73591, 73592, 73593, 73594, 73595, 73596, 73597, 73598, 73599, 73600, 
    73601, 73602, 73603, 73604, 73605, 73606, 73607, 73608, 73609, 73610, 
    73611, 73612, 73613, 73614, 73615, 73616, 73617, 73618, 73619, 73620, 
    73621, 73622, 73623, 73624, 73625, 73626, 73627, 73628, 73629, 73630, 
    73631, 73632, 73633, 73634, 73635, 73636, 73637, 73638, 73639, 73640, 
    73641, 73642, 73643, 73644, 73645, 73646, 73647, 73648, 73649, 73650, 
    73651, 73652, 73653, 73654, 73655, 73656, 73657, 73658, 73659, 73660, 
    73661, 73662, 73663, 73664, 73665, 73666, 73667, 73668, 73669, 73670, 
    73671, 73672, 73673, 73674, 73675, 73676, 73677, 73678, 73679, 73680, 
    73681, 73682, 73683, 73684, 73685, 73686, 73687, 73688, 73689, 73690, 
    73691, 73692, 73693, 73694, 73695, 73696, 73697, 73698, 73699, 73700, 
    73701, 73702, 73703, 73704, 73705, 73706, 73707, 73708, 73709, 73710, 
    73711, 73712, 73713, 73714, 73715, 73716, 73717, 73718, 73719, 73720, 
    73721, 73722, 73723, 73724, 73725, 73726, 73727, 73728, 73729, 73730, 
    73731, 73732, 73733, 73734, 73735, 73736, 73737, 73738, 73739, 73740, 
    73741, 73742, 73743, 73744, 73745, 73746, 73747, 73748, 73749, 73750, 
    73751, 73752, 73753, 73754, 73755, 73756, 73757, 73758, 73759, 73760, 
    73761, 73762, 73763, 73764, 73765, 73766, 73767, 73768, 73769, 73770, 
    73771, 73772, 73773, 73774, 73775, 73776, 73777, 73778, 73779, 73780, 
    73781, 73782, 73783, 73784, 73785, 73786, 73787, 73788, 73789, 73790, 
    73791, 73792, 73793, 73794, 73795, 73796, 73797, 73798, 73799, 73800, 
    73801, 73802, 73803, 73804, 73805, 73806, 73807, 73808, 73809, 73810, 
    73811, 73812, 73813, 73814, 73815, 73816, 73817, 73818, 73819, 73820, 
    73821, 73822, 73823, 73824, 73825, 73826, 73827, 73828, 73829, 73830, 
    73831, 73832, 73833, 73834, 73835, 73836, 73837, 73838, 73839, 73840, 
    73841, 73842, 73843, 73844, 73845, 73846, 73847, 73848, 73849, 73850, 
    73851, 73852, 73853, 73854, 73855, 73856, 73857, 73858, 73859, 73860, 
    73861, 73862, 73863, 73864, 73865, 73866, 73867, 73868, 73869, 73870, 
    73871, 73872, 73873, 73874, 73875, 73876, 73877, 73878, 73879, 73880, 
    73881, 73882, 73883, 73884, 73885, 73886, 73887, 73888, 73889, 73890, 
    73891, 73892, 73893, 73894, 73895, 73896, 73897, 73898, 73899, 73900, 
    73901, 73902, 73903, 73904, 73905, 73906, 73907, 73908, 73909, 73910, 
    73911, 73912, 73913, 73914, 73915, 73916, 73917, 73918, 73919, 73920, 
    73921, 73922, 73923, 73924, 73925, 73926, 73927, 73928, 73929, 73930, 
    73931, 73932, 73933, 73934, 73935, 73936, 73937, 73938, 73939, 73940, 
    73941, 73942, 73943, 73944, 73945, 73946, 73947, 73948, 73949, 73950, 
    73951, 73952, 73953, 73954, 73955, 73956, 73957, 73958, 73959, 73960, 
    73961, 73962, 73963, 73964, 73965, 73966, 73967, 73968, 73969, 73970, 
    73971, 73972, 73973, 73974, 73975, 73976, 73977, 73978, 73979, 73980, 
    73981, 73982, 73983, 73984, 73985, 73986, 73987, 73988, 73989, 73990, 
    73991, 73992, 73993, 73994, 73995, 73996, 73997, 73998, 73999, 74000, 
    74001, 74002, 74003, 74004, 74005, 74006, 74007, 74008, 74009, 74010, 
    74011, 74012, 74013, 74014, 74015, 74016, 74017, 74018, 74019, 74020, 
    74021, 74022, 74023, 74024, 74025, 74026, 74027, 74028, 74029, 74030, 
    74031, 74032, 74033, 74034, 74035, 74036, 74037, 74038, 74039, 74040, 
    74041, 74042, 74043, 74044, 74045, 74046, 74047, 74048, 74049, 74050, 
    74051, 74052, 74053, 74054, 74055, 74056, 74057, 74058, 74059, 74060, 
    74061, 74062, 74063, 74064, 74065, 74066, 74067, 74068, 74069, 74070, 
    74071, 74072, 74073, 74074, 74075, 74076, 74077, 74078, 74079, 74080, 
    74081, 74082, 74083, 74084, 74085, 74086, 74087, 74088, 74089, 74090, 
    74091, 74092, 74093, 74094, 74095, 74096, 74097, 74098, 74099, 74100, 
    74101, 74102, 74103, 74104, 74105, 74106, 74107, 74108, 74109, 74110, 
    74111, 74112, 74113, 74114, 74115, 74116, 74117, 74118, 74119, 74120, 
    74121, 74122, 74123, 74124, 74125, 74126, 74127, 74128, 74129, 74130, 
    74131, 74132, 74133, 74134, 74135, 74136, 74137, 74138, 74139, 74140, 
    74141, 74142, 74143, 74144, 74145, 74146, 74147, 74148, 74149, 74150, 
    74151, 74152, 74153, 74154, 74155, 74156, 74157, 74158, 74159, 74160, 
    74161, 74162, 74163, 74164, 74165, 74166, 74167, 74168, 74169, 74170, 
    74171, 74172, 74173, 74174, 74175, 74176, 74177, 74178, 74179, 74180, 
    74181, 74182, 74183, 74184, 74185, 74186, 74187, 74188, 74189, 74190, 
    74191, 74192, 74193, 74194, 74195, 74196, 74197, 74198, 74199, 74200, 
    74201, 74202, 74203, 74204, 74205, 74206, 74207, 74208, 74209, 74210, 
    74211, 74212, 74213, 74214, 74215, 74216, 74217, 74218, 74219, 74220, 
    74221, 74222, 74223, 74224, 74225, 74226, 74227, 74228, 74229, 74230, 
    74231, 74232, 74233, 74234, 74235, 74236, 74237, 74238, 74239, 74240, 
    74241, 74242, 74243, 74244, 74245, 74246, 74247, 74248, 74249, 74250, 
    74251, 74252, 74253, 74254, 74255, 74256, 74257, 74258, 74259, 74260, 
    74261, 74262, 74263, 74264, 74265, 74266, 74267, 74268, 74269, 74270, 
    74271, 74272, 74273, 74274, 74275, 74276, 74277, 74278, 74279, 74280, 
    74281, 74282, 74283, 74284, 74285, 74286, 74287, 74288, 74289, 74290, 
    74291, 74292, 74293, 74294, 74295, 74296, 74297, 74298, 74299, 74300, 
    74301, 74302, 74303, 74304, 74305, 74306, 74307, 74308, 74309, 74310, 
    74311, 74312, 74313, 74314, 74315, 74316, 74317, 74318, 74319, 74320, 
    74321, 74322, 74323, 74324, 74325, 74326, 74327, 74328, 74329, 74330, 
    74331, 74332, 74333, 74334, 74335, 74336, 74337, 74338, 74339, 74340, 
    74341, 74342, 74343, 74344, 74345, 74346, 74347, 74348, 74349, 74350, 
    74351, 74352, 74353, 74354, 74355, 74356, 74357, 74358, 74359, 74360, 
    74361, 74362, 74363, 74364, 74365, 74366, 74367, 74368, 74369, 74370, 
    74371, 74372, 74373, 74374, 74375, 74376, 74377, 74378, 74379, 74380, 
    74381, 74382, 74383, 74384, 74385, 74386, 74387, 74388, 74389, 74390, 
    74391, 74392, 74393, 74394, 74395, 74396, 74397, 74398, 74399, 74400, 
    74401, 74402, 74403, 74404, 74405, 74406, 74407, 74408, 74409, 74410, 
    74411, 74412, 74413, 74414, 74415, 74416, 74417, 74418, 74419, 74420, 
    74421, 74422, 74423, 74424, 74425, 74426, 74427, 74428, 74429, 74430, 
    74431, 74432, 74433, 74434, 74435, 74436, 74437, 74438, 74439, 74440, 
    74441, 74442, 74443, 74444, 74445, 74446, 74447, 74448, 74449, 74450, 
    74451, 74452, 74453, 74454, 74455, 74456, 74457, 74458, 74459, 74460, 
    74461, 74462, 74463, 74464, 74465, 74466, 74467, 74468, 74469, 74470, 
    74471, 74472, 74473, 74474, 74475, 74476, 74477, 74478, 74479, 74480, 
    74481, 74482, 74483, 74484, 74485, 74486, 74487, 74488, 74489, 74490, 
    74491, 74492, 74493, 74494, 74495, 74496, 74497, 74498, 74499, 74500, 
    74501, 74502, 74503, 74504, 74505, 74506, 74507, 74508, 74509, 74510, 
    74511, 74512, 74513, 74514, 74515, 74516, 74517, 74518, 74519, 74520, 
    74521, 74522, 74523, 74524, 74525, 74526, 74527, 74528, 74529, 74530, 
    74531, 74532, 74533, 74534, 74535, 74536, 74537, 74538, 74539, 74540, 
    74541, 74542, 74543, 74544, 74545, 74546, 74547, 74548, 74549, 74550, 
    74551, 74552, 74553, 74554, 74555, 74556, 74557, 74558, 74559, 74560, 
    74561, 74562, 74563, 74564, 74565, 74566, 74567, 74568, 74569, 74570, 
    74571, 74572, 74573, 74574, 74575, 74576, 74577, 74578, 74579, 74580, 
    74581, 74582, 74583, 74584, 74585, 74586, 74587, 74588, 74589, 74590, 
    74591, 74592, 74593, 74594, 74595, 74596, 74597, 74598, 74599, 74600, 
    74601, 74602, 74603, 74604, 74605, 74606, 74607, 74608, 74609, 74610, 
    74611, 74612, 74613, 74614, 74615, 74616, 74617, 74618, 74619, 74620, 
    74621, 74622, 74623, 74624, 74625, 74626, 74627, 74628, 74629, 74630, 
    74631, 74632, 74633, 74634, 74635, 74636, 74637, 74638, 74639, 74640, 
    74641, 74642, 74643, 74644, 74645, 74646, 74647, 74648, 74649, 74650, 
    74651, 74652, 74653, 74654, 74655, 74656, 74657, 74658, 74659, 74660, 
    74661, 74662, 74663, 74664, 74665, 74666, 74667, 74668, 74669, 74670, 
    74671, 74672, 74673, 74674, 74675, 74676, 74677, 74678, 74679, 74680, 
    74681, 74682, 74683, 74684, 74685, 74686, 74687, 74688, 74689, 74690, 
    74691, 74692, 74693, 74694, 74695, 74696, 74697, 74698, 74699, 74700, 
    74701, 74702, 74703, 74704, 74705, 74706, 74707, 74708, 74709, 74710, 
    74711, 74712, 74713, 74714, 74715, 74716, 74717, 74718, 74719, 74720, 
    74721, 74722, 74723, 74724, 74725, 74726, 74727, 74728, 74729, 74730, 
    74731, 74732, 74733, 74734, 74735, 74736, 74737, 74738, 74739, 74740, 
    74741, 74742, 74743, 74744, 74745, 74746, 74747, 74748, 74749, 74750, 
    74751, 74752, 74753, 74754, 74755, 74756, 74757, 74758, 74759, 74760, 
    74761, 74762, 74763, 74764, 74765, 74766, 74767, 74768, 74769, 74770, 
    74771, 74772, 74773, 74774, 74775, 74776, 74777, 74778, 74779, 74780, 
    74781, 74782, 74783, 74784, 74785, 74786, 74787, 74788, 74789, 74790, 
    74791, 74792, 74793, 74794, 74795, 74796, 74797, 74798, 74799, 74800, 
    74801, 74802, 74803, 74804, 74805, 74806, 74807, 74808, 74809, 74810, 
    74811, 74812, 74813, 74814, 74815, 74816, 74817, 74818, 74819, 74820, 
    74821, 74822, 74823, 74824, 74825, 74826, 74827, 74828, 74829, 74830, 
    74831, 74832, 74833, 74834, 74835, 74836, 74837, 74838, 74839, 74840, 
    74841, 74842, 74843, 74844, 74845, 74846, 74847, 74848, 74849, 74850, 
    74851, 74852, 74853, 74854, 74855, 74856, 74857, 74858, 74859, 74860, 
    74861, 74862, 74863, 74864, 74865, 74866, 74867, 74868, 74869, 74870, 
    74871, 74872, 74873, 74874, 74875, 74876, 74877, 74878, 74879, 74880, 
    74881, 74882, 74883, 74884, 74885, 74886, 74887, 74888, 74889, 74890, 
    74891, 74892, 74893, 74894, 74895, 74896, 74897, 74898, 74899, 74900, 
    74901, 74902, 74903, 74904, 74905, 74906, 74907, 74908, 74909, 74910, 
    74911, 74912, 74913, 74914, 74915, 74916, 74917, 74918, 74919, 74920, 
    74921, 74922, 74923, 74924, 74925, 74926, 74927, 74928, 74929, 74930, 
    74931, 74932, 74933, 74934, 74935, 74936, 74937, 74938, 74939, 74940, 
    74941, 74942, 74943, 74944, 74945, 74946, 74947, 74948, 74949, 74950, 
    74951, 74952, 74953, 74954, 74955, 74956, 74957, 74958, 74959, 74960, 
    74961, 74962, 74963, 74964, 74965, 74966, 74967, 74968, 74969, 74970, 
    74971, 74972, 74973, 74974, 74975, 74976, 74977, 74978, 74979, 74980, 
    74981, 74982, 74983, 74984, 74985, 74986, 74987, 74988, 74989, 74990, 
    74991, 74992, 74993, 74994, 74995, 74996, 74997, 74998, 74999, 75000, 
    75001, 75002, 75003, 75004, 75005, 75006, 75007, 75008, 75009, 75010, 
    75011, 75012, 75013, 75014, 75015, 75016, 75017, 75018, 75019, 75020, 
    75021, 75022, 75023, 75024, 75025, 75026, 75027, 75028, 75029, 75030, 
    75031, 75032, 75033, 75034, 75035, 75036, 75037, 75038, 75039, 75040, 
    75041, 75042, 75043, 75044, 75045, 75046, 75047, 75048, 75049, 75050, 
    75051, 75052, 75053, 75054, 75055, 75056, 75057, 75058, 75059, 75060, 
    75061, 75062, 75063, 75064, 75065, 75066, 75067, 75068, 75069, 75070, 
    75071, 75072, 75073, 75074, 75075, 75076, 75077, 75078, 75079, 75080, 
    75081, 75082, 75083, 75084, 75085, 75086, 75087, 75088, 75089, 75090, 
    75091, 75092, 75093, 75094, 75095, 75096, 75097, 75098, 75099, 75100, 
    75101, 75102, 75103, 75104, 75105, 75106, 75107, 75108, 75109, 75110, 
    75111, 75112, 75113, 75114, 75115, 75116, 75117, 75118, 75119, 75120, 
    75121, 75122, 75123, 75124, 75125, 75126, 75127, 75128, 75129, 75130, 
    75131, 75132, 75133, 75134, 75135, 75136, 75137, 75138, 75139, 75140, 
    75141, 75142, 75143, 75144, 75145, 75146, 75147, 75148, 75149, 75150, 
    75151, 75152, 75153, 75154, 75155, 75156, 75157, 75158, 75159, 75160, 
    75161, 75162, 75163, 75164, 75165, 75166, 75167, 75168, 75169, 75170, 
    75171, 75172, 75173, 75174, 75175, 75176, 75177, 75178, 75179, 75180, 
    75181, 75182, 75183, 75184, 75185, 75186, 75187, 75188, 75189, 75190, 
    75191, 75192, 75193, 75194, 75195, 75196, 75197, 75198, 75199, 75200, 
    75201, 75202, 75203, 75204, 75205, 75206, 75207, 75208, 75209, 75210, 
    75211, 75212, 75213, 75214, 75215, 75216, 75217, 75218, 75219, 75220, 
    75221, 75222, 75223, 75224, 75225, 75226, 75227, 75228, 75229, 75230, 
    75231, 75232, 75233, 75234, 75235, 75236, 75237, 75238, 75239, 75240, 
    75241, 75242, 75243, 75244, 75245, 75246, 75247, 75248, 75249, 75250, 
    75251, 75252, 75253, 75254, 75255, 75256, 75257, 75258, 75259, 75260, 
    75261, 75262, 75263, 75264, 75265, 75266, 75267, 75268, 75269, 75270, 
    75271, 75272, 75273, 75274, 75275, 75276, 75277, 75278, 75279, 75280, 
    75281, 75282, 75283, 75284, 75285, 75286, 75287, 75288, 75289, 75290, 
    75291, 75292, 75293, 75294, 75295, 75296, 75297, 75298, 75299, 75300, 
    75301, 75302, 75303, 75304, 75305, 75306, 75307, 75308, 75309, 75310, 
    75311, 75312, 75313, 75314, 75315, 75316, 75317, 75318, 75319, 75320, 
    75321, 75322, 75323, 75324, 75325, 75326, 75327, 75328, 75329, 75330, 
    75331, 75332, 75333, 75334, 75335, 75336, 75337, 75338, 75339, 75340, 
    75341, 75342, 75343, 75344, 75345, 75346, 75347, 75348, 75349, 75350, 
    75351, 75352, 75353, 75354, 75355, 75356, 75357, 75358, 75359, 75360, 
    75361, 75362, 75363, 75364, 75365, 75366, 75367, 75368, 75369, 75370, 
    75371, 75372, 75373, 75374, 75375, 75376, 75377, 75378, 75379, 75380, 
    75381, 75382, 75383, 75384, 75385, 75386, 75387, 75388, 75389, 75390, 
    75391, 75392, 75393, 75394, 75395, 75396, 75397, 75398, 75399, 75400, 
    75401, 75402, 75403, 75404, 75405, 75406, 75407, 75408, 75409, 75410, 
    75411, 75412, 75413, 75414, 75415, 75416, 75417, 75418, 75419, 75420, 
    75421, 75422, 75423, 75424, 75425, 75426, 75427, 75428, 75429, 75430, 
    75431, 75432, 75433, 75434, 75435, 75436, 75437, 75438, 75439, 75440, 
    75441, 75442, 75443, 75444, 75445, 75446, 75447, 75448, 75449, 75450, 
    75451, 75452, 75453, 75454, 75455, 75456, 75457, 75458, 75459, 75460, 
    75461, 75462, 75463, 75464, 75465, 75466, 75467, 75468, 75469, 75470, 
    75471, 75472, 75473, 75474, 75475, 75476, 75477, 75478, 75479, 75480, 
    75481, 75482, 75483, 75484, 75485, 75486, 75487, 75488, 75489, 75490, 
    75491, 75492, 75493, 75494, 75495, 75496, 75497, 75498, 75499, 75500, 
    75501, 75502, 75503, 75504, 75505, 75506, 75507, 75508, 75509, 75510, 
    75511, 75512, 75513, 75514, 75515, 75516, 75517, 75518, 75519, 75520, 
    75521, 75522, 75523, 75524, 75525, 75526, 75527, 75528, 75529, 75530, 
    75531, 75532, 75533, 75534, 75535, 75536, 75537, 75538, 75539, 75540, 
    75541, 75542, 75543, 75544, 75545, 75546, 75547, 75548, 75549, 75550, 
    75551, 75552, 75553, 75554, 75555, 75556, 75557, 75558, 75559, 75560, 
    75561, 75562, 75563, 75564, 75565, 75566, 75567, 75568, 75569, 75570, 
    75571, 75572, 75573, 75574, 75575, 75576, 75577, 75578, 75579, 75580, 
    75581, 75582, 75583, 75584, 75585, 75586, 75587, 75588, 75589, 75590, 
    75591, 75592, 75593, 75594, 75595, 75596, 75597, 75598, 75599, 75600, 
    75601, 75602, 75603, 75604, 75605, 75606, 75607, 75608, 75609, 75610, 
    75611, 75612, 75613, 75614, 75615, 75616, 75617, 75618, 75619, 75620, 
    75621, 75622, 75623, 75624, 75625, 75626, 75627, 75628, 75629, 75630, 
    75631, 75632, 75633, 75634, 75635, 75636, 75637, 75638, 75639, 75640, 
    75641, 75642, 75643, 75644, 75645, 75646, 75647, 75648, 75649, 75650, 
    75651, 75652, 75653, 75654, 75655, 75656, 75657, 75658, 75659, 75660, 
    75661, 75662, 75663, 75664, 75665, 75666, 75667, 75668, 75669, 75670, 
    75671, 75672, 75673, 75674, 75675, 75676, 75677, 75678, 75679, 75680, 
    75681, 75682, 75683, 75684, 75685, 75686, 75687, 75688, 75689, 75690, 
    75691, 75692, 75693, 75694, 75695, 75696, 75697, 75698, 75699, 75700, 
    75701, 75702, 75703, 75704, 75705, 75706, 75707, 75708, 75709, 75710, 
    75711, 75712, 75713, 75714, 75715, 75716, 75717, 75718, 75719, 75720, 
    75721, 75722, 75723, 75724, 75725, 75726, 75727, 75728, 75729, 75730, 
    75731, 75732, 75733, 75734, 75735, 75736, 75737, 75738, 75739, 75740, 
    75741, 75742, 75743, 75744, 75745, 75746, 75747, 75748, 75749, 75750, 
    75751, 75752, 75753, 75754, 75755, 75756, 75757, 75758, 75759, 75760, 
    75761, 75762, 75763, 75764, 75765, 75766, 75767, 75768, 75769, 75770, 
    75771, 75772, 75773, 75774, 75775, 75776, 75777, 75778, 75779, 75780, 
    75781, 75782, 75783, 75784, 75785, 75786, 75787, 75788, 75789, 75790, 
    75791, 75792, 75793, 75794, 75795, 75796, 75797, 75798, 75799, 75800, 
    75801, 75802, 75803, 75804, 75805, 75806, 75807, 75808, 75809, 75810, 
    75811, 75812, 75813, 75814, 75815, 75816, 75817, 75818, 75819, 75820, 
    75821, 75822, 75823, 75824, 75825, 75826, 75827, 75828, 75829, 75830, 
    75831, 75832, 75833, 75834, 75835, 75836, 75837, 75838, 75839, 75840, 
    75841, 75842, 75843, 75844, 75845, 75846, 75847, 75848, 75849, 75850, 
    75851, 75852, 75853, 75854, 75855, 75856, 75857, 75858, 75859, 75860, 
    75861, 75862, 75863, 75864, 75865, 75866, 75867, 75868, 75869, 75870, 
    75871, 75872, 75873, 75874, 75875, 75876, 75877, 75878, 75879, 75880, 
    75881, 75882, 75883, 75884, 75885, 75886, 75887, 75888, 75889, 75890, 
    75891, 75892, 75893, 75894, 75895, 75896, 75897, 75898, 75899, 75900, 
    75901, 75902, 75903, 75904, 75905, 75906, 75907, 75908, 75909, 75910, 
    75911, 75912, 75913, 75914, 75915, 75916, 75917, 75918, 75919, 75920, 
    75921, 75922, 75923, 75924, 75925, 75926, 75927, 75928, 75929, 75930, 
    75931, 75932, 75933, 75934, 75935, 75936, 75937, 75938, 75939, 75940, 
    75941, 75942, 75943, 75944, 75945, 75946, 75947, 75948, 75949, 75950, 
    75951, 75952, 75953, 75954, 75955, 75956, 75957, 75958, 75959, 75960, 
    75961, 75962, 75963, 75964, 75965, 75966, 75967, 75968, 75969, 75970, 
    75971, 75972, 75973, 75974, 75975, 75976, 75977, 75978, 75979, 75980, 
    75981, 75982, 75983, 75984, 75985, 75986, 75987, 75988, 75989, 75990, 
    75991, 75992, 75993, 75994, 75995, 75996, 75997, 75998, 75999, 76000, 
    76001, 76002, 76003, 76004, 76005, 76006, 76007, 76008, 76009, 76010, 
    76011, 76012, 76013, 76014, 76015, 76016, 76017, 76018, 76019, 76020, 
    76021, 76022, 76023, 76024, 76025, 76026, 76027, 76028, 76029, 76030, 
    76031, 76032, 76033, 76034, 76035, 76036, 76037, 76038, 76039, 76040, 
    76041, 76042, 76043, 76044, 76045, 76046, 76047, 76048, 76049, 76050, 
    76051, 76052, 76053, 76054, 76055, 76056, 76057, 76058, 76059, 76060, 
    76061, 76062, 76063, 76064, 76065, 76066, 76067, 76068, 76069, 76070, 
    76071, 76072, 76073, 76074, 76075, 76076, 76077, 76078, 76079, 76080, 
    76081, 76082, 76083, 76084, 76085, 76086, 76087, 76088, 76089, 76090, 
    76091, 76092, 76093, 76094, 76095, 76096, 76097, 76098, 76099, 76100, 
    76101, 76102, 76103, 76104, 76105, 76106, 76107, 76108, 76109, 76110, 
    76111, 76112, 76113, 76114, 76115, 76116, 76117, 76118, 76119, 76120, 
    76121, 76122, 76123, 76124, 76125, 76126, 76127, 76128, 76129, 76130, 
    76131, 76132, 76133, 76134, 76135, 76136, 76137, 76138, 76139, 76140, 
    76141, 76142, 76143, 76144, 76145, 76146, 76147, 76148, 76149, 76150, 
    76151, 76152, 76153, 76154, 76155, 76156, 76157, 76158, 76159, 76160, 
    76161, 76162, 76163, 76164, 76165, 76166, 76167, 76168, 76169, 76170, 
    76171, 76172, 76173, 76174, 76175, 76176, 76177, 76178, 76179, 76180, 
    76181, 76182, 76183, 76184, 76185, 76186, 76187, 76188, 76189, 76190, 
    76191, 76192, 76193, 76194, 76195, 76196, 76197, 76198, 76199, 76200, 
    76201, 76202, 76203, 76204, 76205, 76206, 76207, 76208, 76209, 76210, 
    76211, 76212, 76213, 76214, 76215, 76216, 76217, 76218, 76219, 76220, 
    76221, 76222, 76223, 76224, 76225, 76226, 76227, 76228, 76229, 76230, 
    76231, 76232, 76233, 76234, 76235, 76236, 76237, 76238, 76239, 76240, 
    76241, 76242, 76243, 76244, 76245, 76246, 76247, 76248, 76249, 76250, 
    76251, 76252, 76253, 76254, 76255, 76256, 76257, 76258, 76259, 76260, 
    76261, 76262, 76263, 76264, 76265, 76266, 76267, 76268, 76269, 76270, 
    76271, 76272, 76273, 76274, 76275, 76276, 76277, 76278, 76279, 76280, 
    76281, 76282, 76283, 76284, 76285, 76286, 76287, 76288, 76289, 76290, 
    76291, 76292, 76293, 76294, 76295, 76296, 76297, 76298, 76299, 76300, 
    76301, 76302, 76303, 76304, 76305, 76306, 76307, 76308, 76309, 76310, 
    76311, 76312, 76313, 76314, 76315, 76316, 76317, 76318, 76319, 76320, 
    76321, 76322, 76323, 76324, 76325, 76326, 76327, 76328, 76329, 76330, 
    76331, 76332, 76333, 76334, 76335, 76336, 76337, 76338, 76339, 76340, 
    76341, 76342, 76343, 76344, 76345, 76346, 76347, 76348, 76349, 76350, 
    76351, 76352, 76353, 76354, 76355, 76356, 76357, 76358, 76359, 76360, 
    76361, 76362, 76363, 76364, 76365, 76366, 76367, 76368, 76369, 76370, 
    76371, 76372, 76373, 76374, 76375, 76376, 76377, 76378, 76379, 76380, 
    76381, 76382, 76383, 76384, 76385, 76386, 76387, 76388, 76389, 76390, 
    76391, 76392, 76393, 76394, 76395, 76396, 76397, 76398, 76399, 76400, 
    76401, 76402, 76403, 76404, 76405, 76406, 76407, 76408, 76409, 76410, 
    76411, 76412, 76413, 76414, 76415, 76416, 76417, 76418, 76419, 76420, 
    76421, 76422, 76423, 76424, 76425, 76426, 76427, 76428, 76429, 76430, 
    76431, 76432, 76433, 76434, 76435, 76436, 76437, 76438, 76439, 76440, 
    76441, 76442, 76443, 76444, 76445, 76446, 76447, 76448, 76449, 76450, 
    76451, 76452, 76453, 76454, 76455, 76456, 76457, 76458, 76459, 76460, 
    76461, 76462, 76463, 76464, 76465, 76466, 76467, 76468, 76469, 76470, 
    76471, 76472, 76473, 76474, 76475, 76476, 76477, 76478, 76479, 76480, 
    76481, 76482, 76483, 76484, 76485, 76486, 76487, 76488, 76489, 76490, 
    76491, 76492, 76493, 76494, 76495, 76496, 76497, 76498, 76499, 76500, 
    76501, 76502, 76503, 76504, 76505, 76506, 76507, 76508, 76509, 76510, 
    76511, 76512, 76513, 76514, 76515, 76516, 76517, 76518, 76519, 76520, 
    76521, 76522, 76523, 76524, 76525, 76526, 76527, 76528, 76529, 76530, 
    76531, 76532, 76533, 76534, 76535, 76536, 76537, 76538, 76539, 76540, 
    76541, 76542, 76543, 76544, 76545, 76546, 76547, 76548, 76549, 76550, 
    76551, 76552, 76553, 76554, 76555, 76556, 76557, 76558, 76559, 76560, 
    76561, 76562, 76563, 76564, 76565, 76566, 76567, 76568, 76569, 76570, 
    76571, 76572, 76573, 76574, 76575, 76576, 76577, 76578, 76579, 76580, 
    76581, 76582, 76583, 76584, 76585, 76586, 76587, 76588, 76589, 76590, 
    76591, 76592, 76593, 76594, 76595, 76596, 76597, 76598, 76599, 76600, 
    76601, 76602, 76603, 76604, 76605, 76606, 76607, 76608, 76609, 76610, 
    76611, 76612, 76613, 76614, 76615, 76616, 76617, 76618, 76619, 76620, 
    76621, 76622, 76623, 76624, 76625, 76626, 76627, 76628, 76629, 76630, 
    76631, 76632, 76633, 76634, 76635, 76636, 76637, 76638, 76639, 76640, 
    76641, 76642, 76643, 76644, 76645, 76646, 76647, 76648, 76649, 76650, 
    76651, 76652, 76653, 76654, 76655, 76656, 76657, 76658, 76659, 76660, 
    76661, 76662, 76663, 76664, 76665, 76666, 76667, 76668, 76669, 76670, 
    76671, 76672, 76673, 76674, 76675, 76676, 76677, 76678, 76679, 76680, 
    76681, 76682, 76683, 76684, 76685, 76686, 76687, 76688, 76689, 76690, 
    76691, 76692, 76693, 76694, 76695, 76696, 76697, 76698, 76699, 76700, 
    76701, 76702, 76703, 76704, 76705, 76706, 76707, 76708, 76709, 76710, 
    76711, 76712, 76713, 76714, 76715, 76716, 76717, 76718, 76719, 76720, 
    76721, 76722, 76723, 76724, 76725, 76726, 76727, 76728, 76729, 76730, 
    76731, 76732, 76733, 76734, 76735, 76736, 76737, 76738, 76739, 76740, 
    76741, 76742, 76743, 76744, 76745, 76746, 76747, 76748, 76749, 76750, 
    76751, 76752, 76753, 76754, 76755, 76756, 76757, 76758, 76759, 76760, 
    76761, 76762, 76763, 76764, 76765, 76766, 76767, 76768, 76769, 76770, 
    76771, 76772, 76773, 76774, 76775, 76776, 76777, 76778, 76779, 76780, 
    76781, 76782, 76783, 76784, 76785, 76786, 76787, 76788, 76789, 76790, 
    76791, 76792, 76793, 76794, 76795, 76796, 76797, 76798, 76799, 76800, 
    76801, 76802, 76803, 76804, 76805, 76806, 76807, 76808, 76809, 76810, 
    76811, 76812, 76813, 76814, 76815, 76816, 76817, 76818, 76819, 76820, 
    76821, 76822, 76823, 76824, 76825, 76826, 76827, 76828, 76829, 76830, 
    76831, 76832, 76833, 76834, 76835, 76836, 76837, 76838, 76839, 76840, 
    76841, 76842, 76843, 76844, 76845, 76846, 76847, 76848, 76849, 76850, 
    76851, 76852, 76853, 76854, 76855, 76856, 76857, 76858, 76859, 76860, 
    76861, 76862, 76863, 76864, 76865, 76866, 76867, 76868, 76869, 76870, 
    76871, 76872, 76873, 76874, 76875, 76876, 76877, 76878, 76879, 76880, 
    76881, 76882, 76883, 76884, 76885, 76886, 76887, 76888, 76889, 76890, 
    76891, 76892, 76893, 76894, 76895, 76896, 76897, 76898, 76899, 76900, 
    76901, 76902, 76903, 76904, 76905, 76906, 76907, 76908, 76909, 76910, 
    76911, 76912, 76913, 76914, 76915, 76916, 76917, 76918, 76919, 76920, 
    76921, 76922, 76923, 76924, 76925, 76926, 76927, 76928, 76929, 76930, 
    76931, 76932, 76933, 76934, 76935, 76936, 76937, 76938, 76939, 76940, 
    76941, 76942, 76943, 76944, 76945, 76946, 76947, 76948, 76949, 76950, 
    76951, 76952, 76953, 76954, 76955, 76956, 76957, 76958, 76959, 76960, 
    76961, 76962, 76963, 76964, 76965, 76966, 76967, 76968, 76969, 76970, 
    76971, 76972, 76973, 76974, 76975, 76976, 76977, 76978, 76979, 76980, 
    76981, 76982, 76983, 76984, 76985, 76986, 76987, 76988, 76989, 76990, 
    76991, 76992, 76993, 76994, 76995, 76996, 76997, 76998, 76999, 77000, 
    77001, 77002, 77003, 77004, 77005, 77006, 77007, 77008, 77009, 77010, 
    77011, 77012, 77013, 77014, 77015, 77016, 77017, 77018, 77019, 77020, 
    77021, 77022, 77023, 77024, 77025, 77026, 77027, 77028, 77029, 77030, 
    77031, 77032, 77033, 77034, 77035, 77036, 77037, 77038, 77039, 77040, 
    77041, 77042, 77043, 77044, 77045, 77046, 77047, 77048, 77049, 77050, 
    77051, 77052, 77053, 77054, 77055, 77056, 77057, 77058, 77059, 77060, 
    77061, 77062, 77063, 77064, 77065, 77066, 77067, 77068, 77069, 77070, 
    77071, 77072, 77073, 77074, 77075, 77076, 77077, 77078, 77079, 77080, 
    77081, 77082, 77083, 77084, 77085, 77086, 77087, 77088, 77089, 77090, 
    77091, 77092, 77093, 77094, 77095, 77096, 77097, 77098, 77099, 77100, 
    77101, 77102, 77103, 77104, 77105, 77106, 77107, 77108, 77109, 77110, 
    77111, 77112, 77113, 77114, 77115, 77116, 77117, 77118, 77119, 77120, 
    77121, 77122, 77123, 77124, 77125, 77126, 77127, 77128, 77129, 77130, 
    77131, 77132, 77133, 77134, 77135, 77136, 77137, 77138, 77139, 77140, 
    77141, 77142, 77143, 77144, 77145, 77146, 77147, 77148, 77149, 77150, 
    77151, 77152, 77153, 77154, 77155, 77156, 77157, 77158, 77159, 77160, 
    77161, 77162, 77163, 77164, 77165, 77166, 77167, 77168, 77169, 77170, 
    77171, 77172, 77173, 77174, 77175, 77176, 77177, 77178, 77179, 77180, 
    77181, 77182, 77183, 77184, 77185, 77186, 77187, 77188, 77189, 77190, 
    77191, 77192, 77193, 77194, 77195, 77196, 77197, 77198, 77199, 77200, 
    77201, 77202, 77203, 77204, 77205, 77206, 77207, 77208, 77209, 77210, 
    77211, 77212, 77213, 77214, 77215, 77216, 77217, 77218, 77219, 77220, 
    77221, 77222, 77223, 77224, 77225, 77226, 77227, 77228, 77229, 77230, 
    77231, 77232, 77233, 77234, 77235, 77236, 77237, 77238, 77239, 77240, 
    77241, 77242, 77243, 77244, 77245, 77246, 77247, 77248, 77249, 77250, 
    77251, 77252, 77253, 77254, 77255, 77256, 77257, 77258, 77259, 77260, 
    77261, 77262, 77263, 77264, 77265, 77266, 77267, 77268, 77269, 77270, 
    77271, 77272, 77273, 77274, 77275, 77276, 77277, 77278, 77279, 77280, 
    77281, 77282, 77283, 77284, 77285, 77286, 77287, 77288, 77289, 77290, 
    77291, 77292, 77293, 77294, 77295, 77296, 77297, 77298, 77299, 77300, 
    77301, 77302, 77303, 77304, 77305, 77306, 77307, 77308, 77309, 77310, 
    77311, 77312, 77313, 77314, 77315, 77316, 77317, 77318, 77319, 77320, 
    77321, 77322, 77323, 77324, 77325, 77326, 77327, 77328, 77329, 77330, 
    77331, 77332, 77333, 77334, 77335, 77336, 77337, 77338, 77339, 77340, 
    77341, 77342, 77343, 77344, 77345, 77346, 77347, 77348, 77349, 77350, 
    77351, 77352, 77353, 77354, 77355, 77356, 77357, 77358, 77359, 77360, 
    77361, 77362, 77363, 77364, 77365, 77366, 77367, 77368, 77369, 77370, 
    77371, 77372, 77373, 77374, 77375, 77376, 77377, 77378, 77379, 77380, 
    77381, 77382, 77383, 77384, 77385, 77386, 77387, 77388, 77389, 77390, 
    77391, 77392, 77393, 77394, 77395, 77396, 77397, 77398, 77399, 77400, 
    77401, 77402, 77403, 77404, 77405, 77406, 77407, 77408, 77409, 77410, 
    77411, 77412, 77413, 77414, 77415, 77416, 77417, 77418, 77419, 77420, 
    77421, 77422, 77423, 77424, 77425, 77426, 77427, 77428, 77429, 77430, 
    77431, 77432, 77433, 77434, 77435, 77436, 77437, 77438, 77439, 77440, 
    77441, 77442, 77443, 77444, 77445, 77446, 77447, 77448, 77449, 77450, 
    77451, 77452, 77453, 77454, 77455, 77456, 77457, 77458, 77459, 77460, 
    77461, 77462, 77463, 77464, 77465, 77466, 77467, 77468, 77469, 77470, 
    77471, 77472, 77473, 77474, 77475, 77476, 77477, 77478, 77479, 77480, 
    77481, 77482, 77483, 77484, 77485, 77486, 77487, 77488, 77489, 77490, 
    77491, 77492, 77493, 77494, 77495, 77496, 77497, 77498, 77499, 77500, 
    77501, 77502, 77503, 77504, 77505, 77506, 77507, 77508, 77509, 77510, 
    77511, 77512, 77513, 77514, 77515, 77516, 77517, 77518, 77519, 77520, 
    77521, 77522, 77523, 77524, 77525, 77526, 77527, 77528, 77529, 77530, 
    77531, 77532, 77533, 77534, 77535, 77536, 77537, 77538, 77539, 77540, 
    77541, 77542, 77543, 77544, 77545, 77546, 77547, 77548, 77549, 77550, 
    77551, 77552, 77553, 77554, 77555, 77556, 77557, 77558, 77559, 77560, 
    77561, 77562, 77563, 77564, 77565, 77566, 77567, 77568, 77569, 77570, 
    77571, 77572, 77573, 77574, 77575, 77576, 77577, 77578, 77579, 77580, 
    77581, 77582, 77583, 77584, 77585, 77586, 77587, 77588, 77589, 77590, 
    77591, 77592, 77593, 77594, 77595, 77596, 77597, 77598, 77599, 77600, 
    77601, 77602, 77603, 77604, 77605, 77606, 77607, 77608, 77609, 77610, 
    77611, 77612, 77613, 77614, 77615, 77616, 77617, 77618, 77619, 77620, 
    77621, 77622, 77623, 77624, 77625, 77626, 77627, 77628, 77629, 77630, 
    77631, 77632, 77633, 77634, 77635, 77636, 77637, 77638, 77639, 77640, 
    77641, 77642, 77643, 77644, 77645, 77646, 77647, 77648, 77649, 77650, 
    77651, 77652, 77653, 77654, 77655, 77656, 77657, 77658, 77659, 77660, 
    77661, 77662, 77663, 77664, 77665, 77666, 77667, 77668, 77669, 77670, 
    77671, 77672, 77673, 77674, 77675, 77676, 77677, 77678, 77679, 77680, 
    77681, 77682, 77683, 77684, 77685, 77686, 77687, 77688, 77689, 77690, 
    77691, 77692, 77693, 77694, 77695, 77696, 77697, 77698, 77699, 77700, 
    77701, 77702, 77703, 77704, 77705, 77706, 77707, 77708, 77709, 77710, 
    77711, 77712, 77713, 77714, 77715, 77716, 77717, 77718, 77719, 77720, 
    77721, 77722, 77723, 77724, 77725, 77726, 77727, 77728, 77729, 77730, 
    77731, 77732, 77733, 77734, 77735, 77736, 77737, 77738, 77739, 77740, 
    77741, 77742, 77743, 77744, 77745, 77746, 77747, 77748, 77749, 77750, 
    77751, 77752, 77753, 77754, 77755, 77756, 77757, 77758, 77759, 77760, 
    77761, 77762, 77763, 77764, 77765, 77766, 77767, 77768, 77769, 77770, 
    77771, 77772, 77773, 77774, 77775, 77776, 77777, 77778, 77779, 77780, 
    77781, 77782, 77783, 77784, 77785, 77786, 77787, 77788, 77789, 77790, 
    77791, 77792, 77793, 77794, 77795, 77796, 77797, 77798, 77799, 77800, 
    77801, 77802, 77803, 77804, 77805, 77806, 77807, 77808, 77809, 77810, 
    77811, 77812, 77813, 77814, 77815, 77816, 77817, 77818, 77819, 77820, 
    77821, 77822, 77823, 77824, 77825, 77826, 77827, 77828, 77829, 77830, 
    77831, 77832, 77833, 77834, 77835, 77836, 77837, 77838, 77839, 77840, 
    77841, 77842, 77843, 77844, 77845, 77846, 77847, 77848, 77849, 77850, 
    77851, 77852, 77853, 77854, 77855, 77856, 77857, 77858, 77859, 77860, 
    77861, 77862, 77863, 77864, 77865, 77866, 77867, 77868, 77869, 77870, 
    77871, 77872, 77873, 77874, 77875, 77876, 77877, 77878, 77879, 77880, 
    77881, 77882, 77883, 77884, 77885, 77886, 77887, 77888, 77889, 77890, 
    77891, 77892, 77893, 77894, 77895, 77896, 77897, 77898, 77899, 77900, 
    77901, 77902, 77903, 77904, 77905, 77906, 77907, 77908, 77909, 77910, 
    77911, 77912, 77913, 77914, 77915, 77916, 77917, 77918, 77919, 77920, 
    77921, 77922, 77923, 77924, 77925, 77926, 77927, 77928, 77929, 77930, 
    77931, 77932, 77933, 77934, 77935, 77936, 77937, 77938, 77939, 77940, 
    77941, 77942, 77943, 77944, 77945, 77946, 77947, 77948, 77949, 77950, 
    77951, 77952, 77953, 77954, 77955, 77956, 77957, 77958, 77959, 77960, 
    77961, 77962, 77963, 77964, 77965, 77966, 77967, 77968, 77969, 77970, 
    77971, 77972, 77973, 77974, 77975, 77976, 77977, 77978, 77979, 77980, 
    77981, 77982, 77983, 77984, 77985, 77986, 77987, 77988, 77989, 77990, 
    77991, 77992, 77993, 77994, 77995, 77996, 77997, 77998, 77999, 78000, 
    78001, 78002, 78003, 78004, 78005, 78006, 78007, 78008, 78009, 78010, 
    78011, 78012, 78013, 78014, 78015, 78016, 78017, 78018, 78019, 78020, 
    78021, 78022, 78023, 78024, 78025, 78026, 78027, 78028, 78029, 78030, 
    78031, 78032, 78033, 78034, 78035, 78036, 78037, 78038, 78039, 78040, 
    78041, 78042, 78043, 78044, 78045, 78046, 78047, 78048, 78049, 78050, 
    78051, 78052, 78053, 78054, 78055, 78056, 78057, 78058, 78059, 78060, 
    78061, 78062, 78063, 78064, 78065, 78066, 78067, 78068, 78069, 78070, 
    78071, 78072, 78073, 78074, 78075, 78076, 78077, 78078, 78079, 78080, 
    78081, 78082, 78083, 78084, 78085, 78086, 78087, 78088, 78089, 78090, 
    78091, 78092, 78093, 78094, 78095, 78096, 78097, 78098, 78099, 78100, 
    78101, 78102, 78103, 78104, 78105, 78106, 78107, 78108, 78109, 78110, 
    78111, 78112, 78113, 78114, 78115, 78116, 78117, 78118, 78119, 78120, 
    78121, 78122, 78123, 78124, 78125, 78126, 78127, 78128, 78129, 78130, 
    78131, 78132, 78133, 78134, 78135, 78136, 78137, 78138, 78139, 78140, 
    78141, 78142, 78143, 78144, 78145, 78146, 78147, 78148, 78149, 78150, 
    78151, 78152, 78153, 78154, 78155, 78156, 78157, 78158, 78159, 78160, 
    78161, 78162, 78163, 78164, 78165, 78166, 78167, 78168, 78169, 78170, 
    78171, 78172, 78173, 78174, 78175, 78176, 78177, 78178, 78179, 78180, 
    78181, 78182, 78183, 78184, 78185, 78186, 78187, 78188, 78189, 78190, 
    78191, 78192, 78193, 78194, 78195, 78196, 78197, 78198, 78199, 78200, 
    78201, 78202, 78203, 78204, 78205, 78206, 78207, 78208, 78209, 78210, 
    78211, 78212, 78213, 78214, 78215, 78216, 78217, 78218, 78219, 78220, 
    78221, 78222, 78223, 78224, 78225, 78226, 78227, 78228, 78229, 78230, 
    78231, 78232, 78233, 78234, 78235, 78236, 78237, 78238, 78239, 78240, 
    78241, 78242, 78243, 78244, 78245, 78246, 78247, 78248, 78249, 78250, 
    78251, 78252, 78253, 78254, 78255, 78256, 78257, 78258, 78259, 78260, 
    78261, 78262, 78263, 78264, 78265, 78266, 78267, 78268, 78269, 78270, 
    78271, 78272, 78273, 78274, 78275, 78276, 78277, 78278, 78279, 78280, 
    78281, 78282, 78283, 78284, 78285, 78286, 78287, 78288, 78289, 78290, 
    78291, 78292, 78293, 78294, 78295, 78296, 78297, 78298, 78299, 78300, 
    78301, 78302, 78303, 78304, 78305, 78306, 78307, 78308, 78309, 78310, 
    78311, 78312, 78313, 78314, 78315, 78316, 78317, 78318, 78319, 78320, 
    78321, 78322, 78323, 78324, 78325, 78326, 78327, 78328, 78329, 78330, 
    78331, 78332, 78333, 78334, 78335, 78336, 78337, 78338, 78339, 78340, 
    78341, 78342, 78343, 78344, 78345, 78346, 78347, 78348, 78349, 78350, 
    78351, 78352, 78353, 78354, 78355, 78356, 78357, 78358, 78359, 78360, 
    78361, 78362, 78363, 78364, 78365, 78366, 78367, 78368, 78369, 78370, 
    78371, 78372, 78373, 78374, 78375, 78376, 78377, 78378, 78379, 78380, 
    78381, 78382, 78383, 78384, 78385, 78386, 78387, 78388, 78389, 78390, 
    78391, 78392, 78393, 78394, 78395, 78396, 78397, 78398, 78399, 78400, 
    78401, 78402, 78403, 78404, 78405, 78406, 78407, 78408, 78409, 78410, 
    78411, 78412, 78413, 78414, 78415, 78416, 78417, 78418, 78419, 78420, 
    78421, 78422, 78423, 78424, 78425, 78426, 78427, 78428, 78429, 78430, 
    78431, 78432, 78433, 78434, 78435, 78436, 78437, 78438, 78439, 78440, 
    78441, 78442, 78443, 78444, 78445, 78446, 78447, 78448, 78449, 78450, 
    78451, 78452, 78453, 78454, 78455, 78456, 78457, 78458, 78459, 78460, 
    78461, 78462, 78463, 78464, 78465, 78466, 78467, 78468, 78469, 78470, 
    78471, 78472, 78473, 78474, 78475, 78476, 78477, 78478, 78479, 78480, 
    78481, 78482, 78483, 78484, 78485, 78486, 78487, 78488, 78489, 78490, 
    78491, 78492, 78493, 78494, 78495, 78496, 78497, 78498, 78499, 78500, 
    78501, 78502, 78503, 78504, 78505, 78506, 78507, 78508, 78509, 78510, 
    78511, 78512, 78513, 78514, 78515, 78516, 78517, 78518, 78519, 78520, 
    78521, 78522, 78523, 78524, 78525, 78526, 78527, 78528, 78529, 78530, 
    78531, 78532, 78533, 78534, 78535, 78536, 78537, 78538, 78539, 78540, 
    78541, 78542, 78543, 78544, 78545, 78546, 78547, 78548, 78549, 78550, 
    78551, 78552, 78553, 78554, 78555, 78556, 78557, 78558, 78559, 78560, 
    78561, 78562, 78563, 78564, 78565, 78566, 78567, 78568, 78569, 78570, 
    78571, 78572, 78573, 78574, 78575, 78576, 78577, 78578, 78579, 78580, 
    78581, 78582, 78583, 78584, 78585, 78586, 78587, 78588, 78589, 78590, 
    78591, 78592, 78593, 78594, 78595, 78596, 78597, 78598, 78599, 78600, 
    78601, 78602, 78603, 78604, 78605, 78606, 78607, 78608, 78609, 78610, 
    78611, 78612, 78613, 78614, 78615, 78616, 78617, 78618, 78619, 78620, 
    78621, 78622, 78623, 78624, 78625, 78626, 78627, 78628, 78629, 78630, 
    78631, 78632, 78633, 78634, 78635, 78636, 78637, 78638, 78639, 78640, 
    78641, 78642, 78643, 78644, 78645, 78646, 78647, 78648, 78649, 78650, 
    78651, 78652, 78653, 78654, 78655, 78656, 78657, 78658, 78659, 78660, 
    78661, 78662, 78663, 78664, 78665, 78666, 78667, 78668, 78669, 78670, 
    78671, 78672, 78673, 78674, 78675, 78676, 78677, 78678, 78679, 78680, 
    78681, 78682, 78683, 78684, 78685, 78686, 78687, 78688, 78689, 78690, 
    78691, 78692, 78693, 78694, 78695, 78696, 78697, 78698, 78699, 78700, 
    78701, 78702, 78703, 78704, 78705, 78706, 78707, 78708, 78709, 78710, 
    78711, 78712, 78713, 78714, 78715, 78716, 78717, 78718, 78719, 78720, 
    78721, 78722, 78723, 78724, 78725, 78726, 78727, 78728, 78729, 78730, 
    78731, 78732, 78733, 78734, 78735, 78736, 78737, 78738, 78739, 78740, 
    78741, 78742, 78743, 78744, 78745, 78746, 78747, 78748, 78749, 78750, 
    78751, 78752, 78753, 78754, 78755, 78756, 78757, 78758, 78759, 78760, 
    78761, 78762, 78763, 78764, 78765, 78766, 78767, 78768, 78769, 78770, 
    78771, 78772, 78773, 78774, 78775, 78776, 78777, 78778, 78779, 78780, 
    78781, 78782, 78783, 78784, 78785, 78786, 78787, 78788, 78789, 78790, 
    78791, 78792, 78793, 78794, 78795, 78796, 78797, 78798, 78799, 78800, 
    78801, 78802, 78803, 78804, 78805, 78806, 78807, 78808, 78809, 78810, 
    78811, 78812, 78813, 78814, 78815, 78816, 78817, 78818, 78819, 78820, 
    78821, 78822, 78823, 78824, 78825, 78826, 78827, 78828, 78829, 78830, 
    78831, 78832, 78833, 78834, 78835, 78836, 78837, 78838, 78839, 78840, 
    78841, 78842, 78843, 78844, 78845, 78846, 78847, 78848, 78849, 78850, 
    78851, 78852, 78853, 78854, 78855, 78856, 78857, 78858, 78859, 78860, 
    78861, 78862, 78863, 78864, 78865, 78866, 78867, 78868, 78869, 78870, 
    78871, 78872, 78873, 78874, 78875, 78876, 78877, 78878, 78879, 78880, 
    78881, 78882, 78883, 78884, 78885, 78886, 78887, 78888, 78889, 78890, 
    78891, 78892, 78893, 78894, 78895, 78896, 78897, 78898, 78899, 78900, 
    78901, 78902, 78903, 78904, 78905, 78906, 78907, 78908, 78909, 78910, 
    78911, 78912, 78913, 78914, 78915, 78916, 78917, 78918, 78919, 78920, 
    78921, 78922, 78923, 78924, 78925, 78926, 78927, 78928, 78929, 78930, 
    78931, 78932, 78933, 78934, 78935, 78936, 78937, 78938, 78939, 78940, 
    78941, 78942, 78943, 78944, 78945, 78946, 78947, 78948, 78949, 78950, 
    78951, 78952, 78953, 78954, 78955, 78956, 78957, 78958, 78959, 78960, 
    78961, 78962, 78963, 78964, 78965, 78966, 78967, 78968, 78969, 78970, 
    78971, 78972, 78973, 78974, 78975, 78976, 78977, 78978, 78979, 78980, 
    78981, 78982, 78983, 78984, 78985, 78986, 78987, 78988, 78989, 78990, 
    78991, 78992, 78993, 78994, 78995, 78996, 78997, 78998, 78999, 79000, 
    79001, 79002, 79003, 79004, 79005, 79006, 79007, 79008, 79009, 79010, 
    79011, 79012, 79013, 79014, 79015, 79016, 79017, 79018, 79019, 79020, 
    79021, 79022, 79023, 79024, 79025, 79026, 79027, 79028, 79029, 79030, 
    79031, 79032, 79033, 79034, 79035, 79036, 79037, 79038, 79039, 79040, 
    79041, 79042, 79043, 79044, 79045, 79046, 79047, 79048, 79049, 79050, 
    79051, 79052, 79053, 79054, 79055, 79056, 79057, 79058, 79059, 79060, 
    79061, 79062, 79063, 79064, 79065, 79066, 79067, 79068, 79069, 79070, 
    79071, 79072, 79073, 79074, 79075, 79076, 79077, 79078, 79079, 79080, 
    79081, 79082, 79083, 79084, 79085, 79086, 79087, 79088, 79089, 79090, 
    79091, 79092, 79093, 79094, 79095, 79096, 79097, 79098, 79099, 79100, 
    79101, 79102, 79103, 79104, 79105, 79106, 79107, 79108, 79109, 79110, 
    79111, 79112, 79113, 79114, 79115, 79116, 79117, 79118, 79119, 79120, 
    79121, 79122, 79123, 79124, 79125, 79126, 79127, 79128, 79129, 79130, 
    79131, 79132, 79133, 79134, 79135, 79136, 79137, 79138, 79139, 79140, 
    79141, 79142, 79143, 79144, 79145, 79146, 79147, 79148, 79149, 79150, 
    79151, 79152, 79153, 79154, 79155, 79156, 79157, 79158, 79159, 79160, 
    79161, 79162, 79163, 79164, 79165, 79166, 79167, 79168, 79169, 79170, 
    79171, 79172, 79173, 79174, 79175, 79176, 79177, 79178, 79179, 79180, 
    79181, 79182, 79183, 79184, 79185, 79186, 79187, 79188, 79189, 79190, 
    79191, 79192, 79193, 79194, 79195, 79196, 79197, 79198, 79199, 79200, 
    79201, 79202, 79203, 79204, 79205, 79206, 79207, 79208, 79209, 79210, 
    79211, 79212, 79213, 79214, 79215, 79216, 79217, 79218, 79219, 79220, 
    79221, 79222, 79223, 79224, 79225, 79226, 79227, 79228, 79229, 79230, 
    79231, 79232, 79233, 79234, 79235, 79236, 79237, 79238, 79239, 79240, 
    79241, 79242, 79243, 79244, 79245, 79246, 79247, 79248, 79249, 79250, 
    79251, 79252, 79253, 79254, 79255, 79256, 79257, 79258, 79259, 79260, 
    79261, 79262, 79263, 79264, 79265, 79266, 79267, 79268, 79269, 79270, 
    79271, 79272, 79273, 79274, 79275, 79276, 79277, 79278, 79279, 79280, 
    79281, 79282, 79283, 79284, 79285, 79286, 79287, 79288, 79289, 79290, 
    79291, 79292, 79293, 79294, 79295, 79296, 79297, 79298, 79299, 79300, 
    79301, 79302, 79303, 79304, 79305, 79306, 79307, 79308, 79309, 79310, 
    79311, 79312, 79313, 79314, 79315, 79316, 79317, 79318, 79319, 79320, 
    79321, 79322, 79323, 79324, 79325, 79326, 79327, 79328, 79329, 79330, 
    79331, 79332, 79333, 79334, 79335, 79336, 79337, 79338, 79339, 79340, 
    79341, 79342, 79343, 79344, 79345, 79346, 79347, 79348, 79349, 79350, 
    79351, 79352, 79353, 79354, 79355, 79356, 79357, 79358, 79359, 79360, 
    79361, 79362, 79363, 79364, 79365, 79366, 79367, 79368, 79369, 79370, 
    79371, 79372, 79373, 79374, 79375, 79376, 79377, 79378, 79379, 79380, 
    79381, 79382, 79383, 79384, 79385, 79386, 79387, 79388, 79389, 79390, 
    79391, 79392, 79393, 79394, 79395, 79396, 79397, 79398, 79399, 79400, 
    79401, 79402, 79403, 79404, 79405, 79406, 79407, 79408, 79409, 79410, 
    79411, 79412, 79413, 79414, 79415, 79416, 79417, 79418, 79419, 79420, 
    79421, 79422, 79423, 79424, 79425, 79426, 79427, 79428, 79429, 79430, 
    79431, 79432, 79433, 79434, 79435, 79436, 79437, 79438, 79439, 79440, 
    79441, 79442, 79443, 79444, 79445, 79446, 79447, 79448, 79449, 79450, 
    79451, 79452, 79453, 79454, 79455, 79456, 79457, 79458, 79459, 79460, 
    79461, 79462, 79463, 79464, 79465, 79466, 79467, 79468, 79469, 79470, 
    79471, 79472, 79473, 79474, 79475, 79476, 79477, 79478, 79479, 79480, 
    79481, 79482, 79483, 79484, 79485, 79486, 79487, 79488, 79489, 79490, 
    79491, 79492, 79493, 79494, 79495, 79496, 79497, 79498, 79499, 79500, 
    79501, 79502, 79503, 79504, 79505, 79506, 79507, 79508, 79509, 79510, 
    79511, 79512, 79513, 79514, 79515, 79516, 79517, 79518, 79519, 79520, 
    79521, 79522, 79523, 79524, 79525, 79526, 79527, 79528, 79529, 79530, 
    79531, 79532, 79533, 79534, 79535, 79536, 79537, 79538, 79539, 79540, 
    79541, 79542, 79543, 79544, 79545, 79546, 79547, 79548, 79549, 79550, 
    79551, 79552, 79553, 79554, 79555, 79556, 79557, 79558, 79559, 79560, 
    79561, 79562, 79563, 79564, 79565, 79566, 79567, 79568, 79569, 79570, 
    79571, 79572, 79573, 79574, 79575, 79576, 79577, 79578, 79579, 79580, 
    79581, 79582, 79583, 79584, 79585, 79586, 79587, 79588, 79589, 79590, 
    79591, 79592, 79593, 79594, 79595, 79596, 79597, 79598, 79599, 79600, 
    79601, 79602, 79603, 79604, 79605, 79606, 79607, 79608, 79609, 79610, 
    79611, 79612, 79613, 79614, 79615, 79616, 79617, 79618, 79619, 79620, 
    79621, 79622, 79623, 79624, 79625, 79626, 79627, 79628, 79629, 79630, 
    79631, 79632, 79633, 79634, 79635, 79636, 79637, 79638, 79639, 79640, 
    79641, 79642, 79643, 79644, 79645, 79646, 79647, 79648, 79649, 79650, 
    79651, 79652, 79653, 79654, 79655, 79656, 79657, 79658, 79659, 79660, 
    79661, 79662, 79663, 79664, 79665, 79666, 79667, 79668, 79669, 79670, 
    79671, 79672, 79673, 79674, 79675, 79676, 79677, 79678, 79679, 79680, 
    79681, 79682, 79683, 79684, 79685, 79686, 79687, 79688, 79689, 79690, 
    79691, 79692, 79693, 79694, 79695, 79696, 79697, 79698, 79699, 79700, 
    79701, 79702, 79703, 79704, 79705, 79706, 79707, 79708, 79709, 79710, 
    79711, 79712, 79713, 79714, 79715, 79716, 79717, 79718, 79719, 79720, 
    79721, 79722, 79723, 79724, 79725, 79726, 79727, 79728, 79729, 79730, 
    79731, 79732, 79733, 79734, 79735, 79736, 79737, 79738, 79739, 79740, 
    79741, 79742, 79743, 79744, 79745, 79746, 79747, 79748, 79749, 79750, 
    79751, 79752, 79753, 79754, 79755, 79756, 79757, 79758, 79759, 79760, 
    79761, 79762, 79763, 79764, 79765, 79766, 79767, 79768, 79769, 79770, 
    79771, 79772, 79773, 79774, 79775, 79776, 79777, 79778, 79779, 79780, 
    79781, 79782, 79783, 79784, 79785, 79786, 79787, 79788, 79789, 79790, 
    79791, 79792, 79793, 79794, 79795, 79796, 79797, 79798, 79799, 79800, 
    79801, 79802, 79803, 79804, 79805, 79806, 79807, 79808, 79809, 79810, 
    79811, 79812, 79813, 79814, 79815, 79816, 79817, 79818, 79819, 79820, 
    79821, 79822, 79823, 79824, 79825, 79826, 79827, 79828, 79829, 79830, 
    79831, 79832, 79833, 79834, 79835, 79836, 79837, 79838, 79839, 79840, 
    79841, 79842, 79843, 79844, 79845, 79846, 79847, 79848, 79849, 79850, 
    79851, 79852, 79853, 79854, 79855, 79856, 79857, 79858, 79859, 79860, 
    79861, 79862, 79863, 79864, 79865, 79866, 79867, 79868, 79869, 79870, 
    79871, 79872, 79873, 79874, 79875, 79876, 79877, 79878, 79879, 79880, 
    79881, 79882, 79883, 79884, 79885, 79886, 79887, 79888, 79889, 79890, 
    79891, 79892, 79893, 79894, 79895, 79896, 79897, 79898, 79899, 79900, 
    79901, 79902, 79903, 79904, 79905, 79906, 79907, 79908, 79909, 79910, 
    79911, 79912, 79913, 79914, 79915, 79916, 79917, 79918, 79919, 79920, 
    79921, 79922, 79923, 79924, 79925, 79926, 79927, 79928, 79929, 79930, 
    79931, 79932, 79933, 79934, 79935, 79936, 79937, 79938, 79939, 79940, 
    79941, 79942, 79943, 79944, 79945, 79946, 79947, 79948, 79949, 79950, 
    79951, 79952, 79953, 79954, 79955, 79956, 79957, 79958, 79959, 79960, 
    79961, 79962, 79963, 79964, 79965, 79966, 79967, 79968, 79969, 79970, 
    79971, 79972, 79973, 79974, 79975, 79976, 79977, 79978, 79979, 79980, 
    79981, 79982, 79983, 79984, 79985, 79986, 79987, 79988, 79989, 79990, 
    79991, 79992, 79993, 79994, 79995, 79996, 79997, 79998, 79999, 80000, 
    80001, 80002, 80003, 80004, 80005, 80006, 80007, 80008, 80009, 80010, 
    80011, 80012, 80013, 80014, 80015, 80016, 80017, 80018, 80019, 80020, 
    80021, 80022, 80023, 80024, 80025, 80026, 80027, 80028, 80029, 80030, 
    80031, 80032, 80033, 80034, 80035, 80036, 80037, 80038, 80039, 80040, 
    80041, 80042, 80043, 80044, 80045, 80046, 80047, 80048, 80049, 80050, 
    80051, 80052, 80053, 80054, 80055, 80056, 80057, 80058, 80059, 80060, 
    80061, 80062, 80063, 80064, 80065, 80066, 80067, 80068, 80069, 80070, 
    80071, 80072, 80073, 80074, 80075, 80076, 80077, 80078, 80079, 80080, 
    80081, 80082, 80083, 80084, 80085, 80086, 80087, 80088, 80089, 80090, 
    80091, 80092, 80093, 80094, 80095, 80096, 80097, 80098, 80099, 80100, 
    80101, 80102, 80103, 80104, 80105, 80106, 80107, 80108, 80109, 80110, 
    80111, 80112, 80113, 80114, 80115, 80116, 80117, 80118, 80119, 80120, 
    80121, 80122, 80123, 80124, 80125, 80126, 80127, 80128, 80129, 80130, 
    80131, 80132, 80133, 80134, 80135, 80136, 80137, 80138, 80139, 80140, 
    80141, 80142, 80143, 80144, 80145, 80146, 80147, 80148, 80149, 80150, 
    80151, 80152, 80153, 80154, 80155, 80156, 80157, 80158, 80159, 80160, 
    80161, 80162, 80163, 80164, 80165, 80166, 80167, 80168, 80169, 80170, 
    80171, 80172, 80173, 80174, 80175, 80176, 80177, 80178, 80179, 80180, 
    80181, 80182, 80183, 80184, 80185, 80186, 80187, 80188, 80189, 80190, 
    80191, 80192, 80193, 80194, 80195, 80196, 80197, 80198, 80199, 80200, 
    80201, 80202, 80203, 80204, 80205, 80206, 80207, 80208, 80209, 80210, 
    80211, 80212, 80213, 80214, 80215, 80216, 80217, 80218, 80219, 80220, 
    80221, 80222, 80223, 80224, 80225, 80226, 80227, 80228, 80229, 80230, 
    80231, 80232, 80233, 80234, 80235, 80236, 80237, 80238, 80239, 80240, 
    80241, 80242, 80243, 80244, 80245, 80246, 80247, 80248, 80249, 80250, 
    80251, 80252, 80253, 80254, 80255, 80256, 80257, 80258, 80259, 80260, 
    80261, 80262, 80263, 80264, 80265, 80266, 80267, 80268, 80269, 80270, 
    80271, 80272, 80273, 80274, 80275, 80276, 80277, 80278, 80279, 80280, 
    80281, 80282, 80283, 80284, 80285, 80286, 80287, 80288, 80289, 80290, 
    80291, 80292, 80293, 80294, 80295, 80296, 80297, 80298, 80299, 80300, 
    80301, 80302, 80303, 80304, 80305, 80306, 80307, 80308, 80309, 80310, 
    80311, 80312, 80313, 80314, 80315, 80316, 80317, 80318, 80319, 80320, 
    80321, 80322, 80323, 80324, 80325, 80326, 80327, 80328, 80329, 80330, 
    80331, 80332, 80333, 80334, 80335, 80336, 80337, 80338, 80339, 80340, 
    80341, 80342, 80343, 80344, 80345, 80346, 80347, 80348, 80349, 80350, 
    80351, 80352, 80353, 80354, 80355, 80356, 80357, 80358, 80359, 80360, 
    80361, 80362, 80363, 80364, 80365, 80366, 80367, 80368, 80369, 80370, 
    80371, 80372, 80373, 80374, 80375, 80376, 80377, 80378, 80379, 80380, 
    80381, 80382, 80383, 80384, 80385, 80386, 80387, 80388, 80389, 80390, 
    80391, 80392, 80393, 80394, 80395, 80396, 80397, 80398, 80399, 80400, 
    80401, 80402, 80403, 80404, 80405, 80406, 80407, 80408, 80409, 80410, 
    80411, 80412, 80413, 80414, 80415, 80416, 80417, 80418, 80419, 80420, 
    80421, 80422, 80423, 80424, 80425, 80426, 80427, 80428, 80429, 80430, 
    80431, 80432, 80433, 80434, 80435, 80436, 80437, 80438, 80439, 80440, 
    80441, 80442, 80443, 80444, 80445, 80446, 80447, 80448, 80449, 80450, 
    80451, 80452, 80453, 80454, 80455, 80456, 80457, 80458, 80459, 80460, 
    80461, 80462, 80463, 80464, 80465, 80466, 80467, 80468, 80469, 80470, 
    80471, 80472, 80473, 80474, 80475, 80476, 80477, 80478, 80479, 80480, 
    80481, 80482, 80483, 80484, 80485, 80486, 80487, 80488, 80489, 80490, 
    80491, 80492, 80493, 80494, 80495, 80496, 80497, 80498, 80499, 80500, 
    80501, 80502, 80503, 80504, 80505, 80506, 80507, 80508, 80509, 80510, 
    80511, 80512, 80513, 80514, 80515, 80516, 80517, 80518, 80519, 80520, 
    80521, 80522, 80523, 80524, 80525, 80526, 80527, 80528, 80529, 80530, 
    80531, 80532, 80533, 80534, 80535, 80536, 80537, 80538, 80539, 80540, 
    80541, 80542, 80543, 80544, 80545, 80546, 80547, 80548, 80549, 80550, 
    80551, 80552, 80553, 80554, 80555, 80556, 80557, 80558, 80559, 80560, 
    80561, 80562, 80563, 80564, 80565, 80566, 80567, 80568, 80569, 80570, 
    80571, 80572, 80573, 80574, 80575, 80576, 80577, 80578, 80579, 80580, 
    80581, 80582, 80583, 80584, 80585, 80586, 80587, 80588, 80589, 80590, 
    80591, 80592, 80593, 80594, 80595, 80596, 80597, 80598, 80599, 80600, 
    80601, 80602, 80603, 80604, 80605, 80606, 80607, 80608, 80609, 80610, 
    80611, 80612, 80613, 80614, 80615, 80616, 80617, 80618, 80619, 80620, 
    80621, 80622, 80623, 80624, 80625, 80626, 80627, 80628, 80629, 80630, 
    80631, 80632, 80633, 80634, 80635, 80636, 80637, 80638, 80639, 80640, 
    80641, 80642, 80643, 80644, 80645, 80646, 80647, 80648, 80649, 80650, 
    80651, 80652, 80653, 80654, 80655, 80656, 80657, 80658, 80659, 80660, 
    80661, 80662, 80663, 80664, 80665, 80666, 80667, 80668, 80669, 80670, 
    80671, 80672, 80673, 80674, 80675, 80676, 80677, 80678, 80679, 80680, 
    80681, 80682, 80683, 80684, 80685, 80686, 80687, 80688, 80689, 80690, 
    80691, 80692, 80693, 80694, 80695, 80696, 80697, 80698, 80699, 80700, 
    80701, 80702, 80703, 80704, 80705, 80706, 80707, 80708, 80709, 80710, 
    80711, 80712, 80713, 80714, 80715, 80716, 80717, 80718, 80719, 80720, 
    80721, 80722, 80723, 80724, 80725, 80726, 80727, 80728, 80729, 80730, 
    80731, 80732, 80733, 80734, 80735, 80736, 80737, 80738, 80739, 80740, 
    80741, 80742, 80743, 80744, 80745, 80746, 80747, 80748, 80749, 80750, 
    80751, 80752, 80753, 80754, 80755, 80756, 80757, 80758, 80759, 80760, 
    80761, 80762, 80763, 80764, 80765, 80766, 80767, 80768, 80769, 80770, 
    80771, 80772, 80773, 80774, 80775, 80776, 80777, 80778, 80779, 80780, 
    80781, 80782, 80783, 80784, 80785, 80786, 80787, 80788, 80789, 80790, 
    80791, 80792, 80793, 80794, 80795, 80796, 80797, 80798, 80799, 80800, 
    80801, 80802, 80803, 80804, 80805, 80806, 80807, 80808, 80809, 80810, 
    80811, 80812, 80813, 80814, 80815, 80816, 80817, 80818, 80819, 80820, 
    80821, 80822, 80823, 80824, 80825, 80826, 80827, 80828, 80829, 80830, 
    80831, 80832, 80833, 80834, 80835, 80836, 80837, 80838, 80839, 80840, 
    80841, 80842, 80843, 80844, 80845, 80846, 80847, 80848, 80849, 80850, 
    80851, 80852, 80853, 80854, 80855, 80856, 80857, 80858, 80859, 80860, 
    80861, 80862, 80863, 80864, 80865, 80866, 80867, 80868, 80869, 80870, 
    80871, 80872, 80873, 80874, 80875, 80876, 80877, 80878, 80879, 80880, 
    80881, 80882, 80883, 80884, 80885, 80886, 80887, 80888, 80889, 80890, 
    80891, 80892, 80893, 80894, 80895, 80896, 80897, 80898, 80899, 80900, 
    80901, 80902, 80903, 80904, 80905, 80906, 80907, 80908, 80909, 80910, 
    80911, 80912, 80913, 80914, 80915, 80916, 80917, 80918, 80919, 80920, 
    80921, 80922, 80923, 80924, 80925, 80926, 80927, 80928, 80929, 80930, 
    80931, 80932, 80933, 80934, 80935, 80936, 80937, 80938, 80939, 80940, 
    80941, 80942, 80943, 80944, 80945, 80946, 80947, 80948, 80949, 80950, 
    80951, 80952, 80953, 80954, 80955, 80956, 80957, 80958, 80959, 80960, 
    80961, 80962, 80963, 80964, 80965, 80966, 80967, 80968, 80969, 80970, 
    80971, 80972, 80973, 80974, 80975, 80976, 80977, 80978, 80979, 80980, 
    80981, 80982, 80983, 80984, 80985, 80986, 80987, 80988, 80989, 80990, 
    80991, 80992, 80993, 80994, 80995, 80996, 80997, 80998, 80999, 81000, 
    81001, 81002, 81003, 81004, 81005, 81006, 81007, 81008, 81009, 81010, 
    81011, 81012, 81013, 81014, 81015, 81016, 81017, 81018, 81019, 81020, 
    81021, 81022, 81023, 81024, 81025, 81026, 81027, 81028, 81029, 81030, 
    81031, 81032, 81033, 81034, 81035, 81036, 81037, 81038, 81039, 81040, 
    81041, 81042, 81043, 81044, 81045, 81046, 81047, 81048, 81049, 81050, 
    81051, 81052, 81053, 81054, 81055, 81056, 81057, 81058, 81059, 81060, 
    81061, 81062, 81063, 81064, 81065, 81066, 81067, 81068, 81069, 81070, 
    81071, 81072, 81073, 81074, 81075, 81076, 81077, 81078, 81079, 81080, 
    81081, 81082, 81083, 81084, 81085, 81086, 81087, 81088, 81089, 81090, 
    81091, 81092, 81093, 81094, 81095, 81096, 81097, 81098, 81099, 81100, 
    81101, 81102, 81103, 81104, 81105, 81106, 81107, 81108, 81109, 81110, 
    81111, 81112, 81113, 81114, 81115, 81116, 81117, 81118, 81119, 81120, 
    81121, 81122, 81123, 81124, 81125, 81126, 81127, 81128, 81129, 81130, 
    81131, 81132, 81133, 81134, 81135, 81136, 81137, 81138, 81139, 81140, 
    81141, 81142, 81143, 81144, 81145, 81146, 81147, 81148, 81149, 81150, 
    81151, 81152, 81153, 81154, 81155, 81156, 81157, 81158, 81159, 81160, 
    81161, 81162, 81163, 81164, 81165, 81166, 81167, 81168, 81169, 81170, 
    81171, 81172, 81173, 81174, 81175, 81176, 81177, 81178, 81179, 81180, 
    81181, 81182, 81183, 81184, 81185, 81186, 81187, 81188, 81189, 81190, 
    81191, 81192, 81193, 81194, 81195, 81196, 81197, 81198, 81199, 81200, 
    81201, 81202, 81203, 81204, 81205, 81206, 81207, 81208, 81209, 81210, 
    81211, 81212, 81213, 81214, 81215, 81216, 81217, 81218, 81219, 81220, 
    81221, 81222, 81223, 81224, 81225, 81226, 81227, 81228, 81229, 81230, 
    81231, 81232, 81233, 81234, 81235, 81236, 81237, 81238, 81239, 81240, 
    81241, 81242, 81243, 81244, 81245, 81246, 81247, 81248, 81249, 81250, 
    81251, 81252, 81253, 81254, 81255, 81256, 81257, 81258, 81259, 81260, 
    81261, 81262, 81263, 81264, 81265, 81266, 81267, 81268, 81269, 81270, 
    81271, 81272, 81273, 81274, 81275, 81276, 81277, 81278, 81279, 81280, 
    81281, 81282, 81283, 81284, 81285, 81286, 81287, 81288, 81289, 81290, 
    81291, 81292, 81293, 81294, 81295, 81296, 81297, 81298, 81299, 81300, 
    81301, 81302, 81303, 81304, 81305, 81306, 81307, 81308, 81309, 81310, 
    81311, 81312, 81313, 81314, 81315, 81316, 81317, 81318, 81319, 81320, 
    81321, 81322, 81323, 81324, 81325, 81326, 81327, 81328, 81329, 81330, 
    81331, 81332, 81333, 81334, 81335, 81336, 81337, 81338, 81339, 81340, 
    81341, 81342, 81343, 81344, 81345, 81346, 81347, 81348, 81349, 81350, 
    81351, 81352, 81353, 81354, 81355, 81356, 81357, 81358, 81359, 81360, 
    81361, 81362, 81363, 81364, 81365, 81366, 81367, 81368, 81369, 81370, 
    81371, 81372, 81373, 81374, 81375, 81376, 81377, 81378, 81379, 81380, 
    81381, 81382, 81383, 81384, 81385, 81386, 81387, 81388, 81389, 81390, 
    81391, 81392, 81393, 81394, 81395, 81396, 81397, 81398, 81399, 81400, 
    81401, 81402, 81403, 81404, 81405, 81406, 81407, 81408, 81409, 81410, 
    81411, 81412, 81413, 81414, 81415, 81416, 81417, 81418, 81419, 81420, 
    81421, 81422, 81423, 81424, 81425, 81426, 81427, 81428, 81429, 81430, 
    81431, 81432, 81433, 81434, 81435, 81436, 81437, 81438, 81439, 81440, 
    81441, 81442, 81443, 81444, 81445, 81446, 81447, 81448, 81449, 81450, 
    81451, 81452, 81453, 81454, 81455, 81456, 81457, 81458, 81459, 81460, 
    81461, 81462, 81463, 81464, 81465, 81466, 81467, 81468, 81469, 81470, 
    81471, 81472, 81473, 81474, 81475, 81476, 81477, 81478, 81479, 81480, 
    81481, 81482, 81483, 81484, 81485, 81486, 81487, 81488, 81489, 81490, 
    81491, 81492, 81493, 81494, 81495, 81496, 81497, 81498, 81499, 81500, 
    81501, 81502, 81503, 81504, 81505, 81506, 81507, 81508, 81509, 81510, 
    81511, 81512, 81513, 81514, 81515, 81516, 81517, 81518, 81519, 81520, 
    81521, 81522, 81523, 81524, 81525, 81526, 81527, 81528, 81529, 81530, 
    81531, 81532, 81533, 81534, 81535, 81536, 81537, 81538, 81539, 81540, 
    81541, 81542, 81543, 81544, 81545, 81546, 81547, 81548, 81549, 81550, 
    81551, 81552, 81553, 81554, 81555, 81556, 81557, 81558, 81559, 81560, 
    81561, 81562, 81563, 81564, 81565, 81566, 81567, 81568, 81569, 81570, 
    81571, 81572, 81573, 81574, 81575, 81576, 81577, 81578, 81579, 81580, 
    81581, 81582, 81583, 81584, 81585, 81586, 81587, 81588, 81589, 81590, 
    81591, 81592, 81593, 81594, 81595, 81596, 81597, 81598, 81599, 81600, 
    81601, 81602, 81603, 81604, 81605, 81606, 81607, 81608, 81609, 81610, 
    81611, 81612, 81613, 81614, 81615, 81616, 81617, 81618, 81619, 81620, 
    81621, 81622, 81623, 81624, 81625, 81626, 81627, 81628, 81629, 81630, 
    81631, 81632, 81633, 81634, 81635, 81636, 81637, 81638, 81639, 81640, 
    81641, 81642, 81643, 81644, 81645, 81646, 81647, 81648, 81649, 81650, 
    81651, 81652, 81653, 81654, 81655, 81656, 81657, 81658, 81659, 81660, 
    81661, 81662, 81663, 81664, 81665, 81666, 81667, 81668, 81669, 81670, 
    81671, 81672, 81673, 81674, 81675, 81676, 81677, 81678, 81679, 81680, 
    81681, 81682, 81683, 81684, 81685, 81686, 81687, 81688, 81689, 81690, 
    81691, 81692, 81693, 81694, 81695, 81696, 81697, 81698, 81699, 81700, 
    81701, 81702, 81703, 81704, 81705, 81706, 81707, 81708, 81709, 81710, 
    81711, 81712, 81713, 81714, 81715, 81716, 81717, 81718, 81719, 81720, 
    81721, 81722, 81723, 81724, 81725, 81726, 81727, 81728, 81729, 81730, 
    81731, 81732, 81733, 81734, 81735, 81736, 81737, 81738, 81739, 81740, 
    81741, 81742, 81743, 81744, 81745, 81746, 81747, 81748, 81749, 81750, 
    81751, 81752, 81753, 81754, 81755, 81756, 81757, 81758, 81759, 81760, 
    81761, 81762, 81763, 81764, 81765, 81766, 81767, 81768, 81769, 81770, 
    81771, 81772, 81773, 81774, 81775, 81776, 81777, 81778, 81779, 81780, 
    81781, 81782, 81783, 81784, 81785, 81786, 81787, 81788, 81789, 81790, 
    81791, 81792, 81793, 81794, 81795, 81796, 81797, 81798, 81799, 81800, 
    81801, 81802, 81803, 81804, 81805, 81806, 81807, 81808, 81809, 81810, 
    81811, 81812, 81813, 81814, 81815, 81816, 81817, 81818, 81819, 81820, 
    81821, 81822, 81823, 81824, 81825, 81826, 81827, 81828, 81829, 81830, 
    81831, 81832, 81833, 81834, 81835, 81836, 81837, 81838, 81839, 81840, 
    81841, 81842, 81843, 81844, 81845, 81846, 81847, 81848, 81849, 81850, 
    81851, 81852, 81853, 81854, 81855, 81856, 81857, 81858, 81859, 81860, 
    81861, 81862, 81863, 81864, 81865, 81866, 81867, 81868, 81869, 81870, 
    81871, 81872, 81873, 81874, 81875, 81876, 81877, 81878, 81879, 81880, 
    81881, 81882, 81883, 81884, 81885, 81886, 81887, 81888, 81889, 81890, 
    81891, 81892, 81893, 81894, 81895, 81896, 81897, 81898, 81899, 81900, 
    81901, 81902, 81903, 81904, 81905, 81906, 81907, 81908, 81909, 81910, 
    81911, 81912, 81913, 81914, 81915, 81916, 81917, 81918, 81919, 81920, 
    81921, 81922, 81923, 81924, 81925, 81926, 81927, 81928, 81929, 81930, 
    81931, 81932, 81933, 81934, 81935, 81936, 81937, 81938, 81939, 81940, 
    81941, 81942, 81943, 81944, 81945, 81946, 81947, 81948, 81949, 81950, 
    81951, 81952, 81953, 81954, 81955, 81956, 81957, 81958, 81959, 81960, 
    81961, 81962, 81963, 81964, 81965, 81966, 81967, 81968, 81969, 81970, 
    81971, 81972, 81973, 81974, 81975, 81976, 81977, 81978, 81979, 81980, 
    81981, 81982, 81983, 81984, 81985, 81986, 81987, 81988, 81989, 81990, 
    81991, 81992, 81993, 81994, 81995, 81996, 81997, 81998, 81999, 82000, 
    82001, 82002, 82003, 82004, 82005, 82006, 82007, 82008, 82009, 82010, 
    82011, 82012, 82013, 82014, 82015, 82016, 82017, 82018, 82019, 82020, 
    82021, 82022, 82023, 82024, 82025, 82026, 82027, 82028, 82029, 82030, 
    82031, 82032, 82033, 82034, 82035, 82036, 82037, 82038, 82039, 82040, 
    82041, 82042, 82043, 82044, 82045, 82046, 82047, 82048, 82049, 82050, 
    82051, 82052, 82053, 82054, 82055, 82056, 82057, 82058, 82059, 82060, 
    82061, 82062, 82063, 82064, 82065, 82066, 82067, 82068, 82069, 82070, 
    82071, 82072, 82073, 82074, 82075, 82076, 82077, 82078, 82079, 82080, 
    82081, 82082, 82083, 82084, 82085, 82086, 82087, 82088, 82089, 82090, 
    82091, 82092, 82093, 82094, 82095, 82096, 82097, 82098, 82099, 82100, 
    82101, 82102, 82103, 82104, 82105, 82106, 82107, 82108, 82109, 82110, 
    82111, 82112, 82113, 82114, 82115, 82116, 82117, 82118, 82119, 82120, 
    82121, 82122, 82123, 82124, 82125, 82126, 82127, 82128, 82129, 82130, 
    82131, 82132, 82133, 82134, 82135, 82136, 82137, 82138, 82139, 82140, 
    82141, 82142, 82143, 82144, 82145, 82146, 82147, 82148, 82149, 82150, 
    82151, 82152, 82153, 82154, 82155, 82156, 82157, 82158, 82159, 82160, 
    82161, 82162, 82163, 82164, 82165, 82166, 82167, 82168, 82169, 82170, 
    82171, 82172, 82173, 82174, 82175, 82176, 82177, 82178, 82179, 82180, 
    82181, 82182, 82183, 82184, 82185, 82186, 82187, 82188, 82189, 82190, 
    82191, 82192, 82193, 82194, 82195, 82196, 82197, 82198, 82199, 82200, 
    82201, 82202, 82203, 82204, 82205, 82206, 82207, 82208, 82209, 82210, 
    82211, 82212, 82213, 82214, 82215, 82216, 82217, 82218, 82219, 82220, 
    82221, 82222, 82223, 82224, 82225, 82226, 82227, 82228, 82229, 82230, 
    82231, 82232, 82233, 82234, 82235, 82236, 82237, 82238, 82239, 82240, 
    82241, 82242, 82243, 82244, 82245, 82246, 82247, 82248, 82249, 82250, 
    82251, 82252, 82253, 82254, 82255, 82256, 82257, 82258, 82259, 82260, 
    82261, 82262, 82263, 82264, 82265, 82266, 82267, 82268, 82269, 82270, 
    82271, 82272, 82273, 82274, 82275, 82276, 82277, 82278, 82279, 82280, 
    82281, 82282, 82283, 82284, 82285, 82286, 82287, 82288, 82289, 82290, 
    82291, 82292, 82293, 82294, 82295, 82296, 82297, 82298, 82299, 82300, 
    82301, 82302, 82303, 82304, 82305, 82306, 82307, 82308, 82309, 82310, 
    82311, 82312, 82313, 82314, 82315, 82316, 82317, 82318, 82319, 82320, 
    82321, 82322, 82323, 82324, 82325, 82326, 82327, 82328, 82329, 82330, 
    82331, 82332, 82333, 82334, 82335, 82336, 82337, 82338, 82339, 82340, 
    82341, 82342, 82343, 82344, 82345, 82346, 82347, 82348, 82349, 82350, 
    82351, 82352, 82353, 82354, 82355, 82356, 82357, 82358, 82359, 82360, 
    82361, 82362, 82363, 82364, 82365, 82366, 82367, 82368, 82369, 82370, 
    82371, 82372, 82373, 82374, 82375, 82376, 82377, 82378, 82379, 82380, 
    82381, 82382, 82383, 82384, 82385, 82386, 82387, 82388, 82389, 82390, 
    82391, 82392, 82393, 82394, 82395, 82396, 82397, 82398, 82399, 82400, 
    82401, 82402, 82403, 82404, 82405, 82406, 82407, 82408, 82409, 82410, 
    82411, 82412, 82413, 82414, 82415, 82416, 82417, 82418, 82419, 82420, 
    82421, 82422, 82423, 82424, 82425, 82426, 82427, 82428, 82429, 82430, 
    82431, 82432, 82433, 82434, 82435, 82436, 82437, 82438, 82439, 82440, 
    82441, 82442, 82443, 82444, 82445, 82446, 82447, 82448, 82449, 82450, 
    82451, 82452, 82453, 82454, 82455, 82456, 82457, 82458, 82459, 82460, 
    82461, 82462, 82463, 82464, 82465, 82466, 82467, 82468, 82469, 82470, 
    82471, 82472, 82473, 82474, 82475, 82476, 82477, 82478, 82479, 82480, 
    82481, 82482, 82483, 82484, 82485, 82486, 82487, 82488, 82489, 82490, 
    82491, 82492, 82493, 82494, 82495, 82496, 82497, 82498, 82499, 82500, 
    82501, 82502, 82503, 82504, 82505, 82506, 82507, 82508, 82509, 82510, 
    82511, 82512, 82513, 82514, 82515, 82516, 82517, 82518, 82519, 82520, 
    82521, 82522, 82523, 82524, 82525, 82526, 82527, 82528, 82529, 82530, 
    82531, 82532, 82533, 82534, 82535, 82536, 82537, 82538, 82539, 82540, 
    82541, 82542, 82543, 82544, 82545, 82546, 82547, 82548, 82549, 82550, 
    82551, 82552, 82553, 82554, 82555, 82556, 82557, 82558, 82559, 82560, 
    82561, 82562, 82563, 82564, 82565, 82566, 82567, 82568, 82569, 82570, 
    82571, 82572, 82573, 82574, 82575, 82576, 82577, 82578, 82579, 82580, 
    82581, 82582, 82583, 82584, 82585, 82586, 82587, 82588, 82589, 82590, 
    82591, 82592, 82593, 82594, 82595, 82596, 82597, 82598, 82599, 82600, 
    82601, 82602, 82603, 82604, 82605, 82606, 82607, 82608, 82609, 82610, 
    82611, 82612, 82613, 82614, 82615, 82616, 82617, 82618, 82619, 82620, 
    82621, 82622, 82623, 82624, 82625, 82626, 82627, 82628, 82629, 82630, 
    82631, 82632, 82633, 82634, 82635, 82636, 82637, 82638, 82639, 82640, 
    82641, 82642, 82643, 82644, 82645, 82646, 82647, 82648, 82649, 82650, 
    82651, 82652, 82653, 82654, 82655, 82656, 82657, 82658, 82659, 82660, 
    82661, 82662, 82663, 82664, 82665, 82666, 82667, 82668, 82669, 82670, 
    82671, 82672, 82673, 82674, 82675, 82676, 82677, 82678, 82679, 82680, 
    82681, 82682, 82683, 82684, 82685, 82686, 82687, 82688, 82689, 82690, 
    82691, 82692, 82693, 82694, 82695, 82696, 82697, 82698, 82699, 82700, 
    82701, 82702, 82703, 82704, 82705, 82706, 82707, 82708, 82709, 82710, 
    82711, 82712, 82713, 82714, 82715, 82716, 82717, 82718, 82719, 82720, 
    82721, 82722, 82723, 82724, 82725, 82726, 82727, 82728, 82729, 82730, 
    82731, 82732, 82733, 82734, 82735, 82736, 82737, 82738, 82739, 82740, 
    82741, 82742, 82743, 82744, 82745, 82746, 82747, 82748, 82749, 82750, 
    82751, 82752, 82753, 82754, 82755, 82756, 82757, 82758, 82759, 82760, 
    82761, 82762, 82763, 82764, 82765, 82766, 82767, 82768, 82769, 82770, 
    82771, 82772, 82773, 82774, 82775, 82776, 82777, 82778, 82779, 82780, 
    82781, 82782, 82783, 82784, 82785, 82786, 82787, 82788, 82789, 82790, 
    82791, 82792, 82793, 82794, 82795, 82796, 82797, 82798, 82799, 82800, 
    82801, 82802, 82803, 82804, 82805, 82806, 82807, 82808, 82809, 82810, 
    82811, 82812, 82813, 82814, 82815, 82816, 82817, 82818, 82819, 82820, 
    82821, 82822, 82823, 82824, 82825, 82826, 82827, 82828, 82829, 82830, 
    82831, 82832, 82833, 82834, 82835, 82836, 82837, 82838, 82839, 82840, 
    82841, 82842, 82843, 82844, 82845, 82846, 82847, 82848, 82849, 82850, 
    82851, 82852, 82853, 82854, 82855, 82856, 82857, 82858, 82859, 82860, 
    82861, 82862, 82863, 82864, 82865, 82866, 82867, 82868, 82869, 82870, 
    82871, 82872, 82873, 82874, 82875, 82876, 82877, 82878, 82879, 82880, 
    82881, 82882, 82883, 82884, 82885, 82886, 82887, 82888, 82889, 82890, 
    82891, 82892, 82893, 82894, 82895, 82896, 82897, 82898, 82899, 82900, 
    82901, 82902, 82903, 82904, 82905, 82906, 82907, 82908, 82909, 82910, 
    82911, 82912, 82913, 82914, 82915, 82916, 82917, 82918, 82919, 82920, 
    82921, 82922, 82923, 82924, 82925, 82926, 82927, 82928, 82929, 82930, 
    82931, 82932, 82933, 82934, 82935, 82936, 82937, 82938, 82939, 82940, 
    82941, 82942, 82943, 82944, 82945, 82946, 82947, 82948, 82949, 82950, 
    82951, 82952, 82953, 82954, 82955, 82956, 82957, 82958, 82959, 82960, 
    82961, 82962, 82963, 82964, 82965, 82966, 82967, 82968, 82969, 82970, 
    82971, 82972, 82973, 82974, 82975, 82976, 82977, 82978, 82979, 82980, 
    82981, 82982, 82983, 82984, 82985, 82986, 82987, 82988, 82989, 82990, 
    82991, 82992, 82993, 82994, 82995, 82996, 82997, 82998, 82999, 83000, 
    83001, 83002, 83003, 83004, 83005, 83006, 83007, 83008, 83009, 83010, 
    83011, 83012, 83013, 83014, 83015, 83016, 83017, 83018, 83019, 83020, 
    83021, 83022, 83023, 83024, 83025, 83026, 83027, 83028, 83029, 83030, 
    83031, 83032, 83033, 83034, 83035, 83036, 83037, 83038, 83039, 83040, 
    83041, 83042, 83043, 83044, 83045, 83046, 83047, 83048, 83049, 83050, 
    83051, 83052, 83053, 83054, 83055, 83056, 83057, 83058, 83059, 83060, 
    83061, 83062, 83063, 83064, 83065, 83066, 83067, 83068, 83069, 83070, 
    83071, 83072, 83073, 83074, 83075, 83076, 83077, 83078, 83079, 83080, 
    83081, 83082, 83083, 83084, 83085, 83086, 83087, 83088, 83089, 83090, 
    83091, 83092, 83093, 83094, 83095, 83096, 83097, 83098, 83099, 83100, 
    83101, 83102, 83103, 83104, 83105, 83106, 83107, 83108, 83109, 83110, 
    83111, 83112, 83113, 83114, 83115, 83116, 83117, 83118, 83119, 83120, 
    83121, 83122, 83123, 83124, 83125, 83126, 83127, 83128, 83129, 83130, 
    83131, 83132, 83133, 83134, 83135, 83136, 83137, 83138, 83139, 83140, 
    83141, 83142, 83143, 83144, 83145, 83146, 83147, 83148, 83149, 83150, 
    83151, 83152, 83153, 83154, 83155, 83156, 83157, 83158, 83159, 83160, 
    83161, 83162, 83163, 83164, 83165, 83166, 83167, 83168, 83169, 83170, 
    83171, 83172, 83173, 83174, 83175, 83176, 83177, 83178, 83179, 83180, 
    83181, 83182, 83183, 83184, 83185, 83186, 83187, 83188, 83189, 83190, 
    83191, 83192, 83193, 83194, 83195, 83196, 83197, 83198, 83199, 83200, 
    83201, 83202, 83203, 83204, 83205, 83206, 83207, 83208, 83209, 83210, 
    83211, 83212, 83213, 83214, 83215, 83216, 83217, 83218, 83219, 83220, 
    83221, 83222, 83223, 83224, 83225, 83226, 83227, 83228, 83229, 83230, 
    83231, 83232, 83233, 83234, 83235, 83236, 83237, 83238, 83239, 83240, 
    83241, 83242, 83243, 83244, 83245, 83246, 83247, 83248, 83249, 83250, 
    83251, 83252, 83253, 83254, 83255, 83256, 83257, 83258, 83259, 83260, 
    83261, 83262, 83263, 83264, 83265, 83266, 83267, 83268, 83269, 83270, 
    83271, 83272, 83273, 83274, 83275, 83276, 83277, 83278, 83279, 83280, 
    83281, 83282, 83283, 83284, 83285, 83286, 83287, 83288, 83289, 83290, 
    83291, 83292, 83293, 83294, 83295, 83296, 83297, 83298, 83299, 83300, 
    83301, 83302, 83303, 83304, 83305, 83306, 83307, 83308, 83309, 83310, 
    83311, 83312, 83313, 83314, 83315, 83316, 83317, 83318, 83319, 83320, 
    83321, 83322, 83323, 83324, 83325, 83326, 83327, 83328, 83329, 83330, 
    83331, 83332, 83333, 83334, 83335, 83336, 83337, 83338, 83339, 83340, 
    83341, 83342, 83343, 83344, 83345, 83346, 83347, 83348, 83349, 83350, 
    83351, 83352, 83353, 83354, 83355, 83356, 83357, 83358, 83359, 83360, 
    83361, 83362, 83363, 83364, 83365, 83366, 83367, 83368, 83369, 83370, 
    83371, 83372, 83373, 83374, 83375, 83376, 83377, 83378, 83379, 83380, 
    83381, 83382, 83383, 83384, 83385, 83386, 83387, 83388, 83389, 83390, 
    83391, 83392, 83393, 83394, 83395, 83396, 83397, 83398, 83399, 83400, 
    83401, 83402, 83403, 83404, 83405, 83406, 83407, 83408, 83409, 83410, 
    83411, 83412, 83413, 83414, 83415, 83416, 83417, 83418, 83419, 83420, 
    83421, 83422, 83423, 83424, 83425, 83426, 83427, 83428, 83429, 83430, 
    83431, 83432, 83433, 83434, 83435, 83436, 83437, 83438, 83439, 83440, 
    83441, 83442, 83443, 83444, 83445, 83446, 83447, 83448, 83449, 83450, 
    83451, 83452, 83453, 83454, 83455, 83456, 83457, 83458, 83459, 83460, 
    83461, 83462, 83463, 83464, 83465, 83466, 83467, 83468, 83469, 83470, 
    83471, 83472, 83473, 83474, 83475, 83476, 83477, 83478, 83479, 83480, 
    83481, 83482, 83483, 83484, 83485, 83486, 83487, 83488, 83489, 83490, 
    83491, 83492, 83493, 83494, 83495, 83496, 83497, 83498, 83499, 83500, 
    83501, 83502, 83503, 83504, 83505, 83506, 83507, 83508, 83509, 83510, 
    83511, 83512, 83513, 83514, 83515, 83516, 83517, 83518, 83519, 83520, 
    83521, 83522, 83523, 83524, 83525, 83526, 83527, 83528, 83529, 83530, 
    83531, 83532, 83533, 83534, 83535, 83536, 83537, 83538, 83539, 83540, 
    83541, 83542, 83543, 83544, 83545, 83546, 83547, 83548, 83549, 83550, 
    83551, 83552, 83553, 83554, 83555, 83556, 83557, 83558, 83559, 83560, 
    83561, 83562, 83563, 83564, 83565, 83566, 83567, 83568, 83569, 83570, 
    83571, 83572, 83573, 83574, 83575, 83576, 83577, 83578, 83579, 83580, 
    83581, 83582, 83583, 83584, 83585, 83586, 83587, 83588, 83589, 83590, 
    83591, 83592, 83593, 83594, 83595, 83596, 83597, 83598, 83599, 83600, 
    83601, 83602, 83603, 83604, 83605, 83606, 83607, 83608, 83609, 83610, 
    83611, 83612, 83613, 83614, 83615, 83616, 83617, 83618, 83619, 83620, 
    83621, 83622, 83623, 83624, 83625, 83626, 83627, 83628, 83629, 83630, 
    83631, 83632, 83633, 83634, 83635, 83636, 83637, 83638, 83639, 83640, 
    83641, 83642, 83643, 83644, 83645, 83646, 83647, 83648, 83649, 83650, 
    83651, 83652, 83653, 83654, 83655, 83656, 83657, 83658, 83659, 83660, 
    83661, 83662, 83663, 83664, 83665, 83666, 83667, 83668, 83669, 83670, 
    83671, 83672, 83673, 83674, 83675, 83676, 83677, 83678, 83679, 83680, 
    83681, 83682, 83683, 83684, 83685, 83686, 83687, 83688, 83689, 83690, 
    83691, 83692, 83693, 83694, 83695, 83696, 83697, 83698, 83699, 83700, 
    83701, 83702, 83703, 83704, 83705, 83706, 83707, 83708, 83709, 83710, 
    83711, 83712, 83713, 83714, 83715, 83716, 83717, 83718, 83719, 83720, 
    83721, 83722, 83723, 83724, 83725, 83726, 83727, 83728, 83729, 83730, 
    83731, 83732, 83733, 83734, 83735, 83736, 83737, 83738, 83739, 83740, 
    83741, 83742, 83743, 83744, 83745, 83746, 83747, 83748, 83749, 83750, 
    83751, 83752, 83753, 83754, 83755, 83756, 83757, 83758, 83759, 83760, 
    83761, 83762, 83763, 83764, 83765, 83766, 83767, 83768, 83769, 83770, 
    83771, 83772, 83773, 83774, 83775, 83776, 83777, 83778, 83779, 83780, 
    83781, 83782, 83783, 83784, 83785, 83786, 83787, 83788, 83789, 83790, 
    83791, 83792, 83793, 83794, 83795, 83796, 83797, 83798, 83799, 83800, 
    83801, 83802, 83803, 83804, 83805, 83806, 83807, 83808, 83809, 83810, 
    83811, 83812, 83813, 83814, 83815, 83816, 83817, 83818, 83819, 83820, 
    83821, 83822, 83823, 83824, 83825, 83826, 83827, 83828, 83829, 83830, 
    83831, 83832, 83833, 83834, 83835, 83836, 83837, 83838, 83839, 83840, 
    83841, 83842, 83843, 83844, 83845, 83846, 83847, 83848, 83849, 83850, 
    83851, 83852, 83853, 83854, 83855, 83856, 83857, 83858, 83859, 83860, 
    83861, 83862, 83863, 83864, 83865, 83866, 83867, 83868, 83869, 83870, 
    83871, 83872, 83873, 83874, 83875, 83876, 83877, 83878, 83879, 83880, 
    83881, 83882, 83883, 83884, 83885, 83886, 83887, 83888, 83889, 83890, 
    83891, 83892, 83893, 83894, 83895, 83896, 83897, 83898, 83899, 83900, 
    83901, 83902, 83903, 83904, 83905, 83906, 83907, 83908, 83909, 83910, 
    83911, 83912, 83913, 83914, 83915, 83916, 83917, 83918, 83919, 83920, 
    83921, 83922, 83923, 83924, 83925, 83926, 83927, 83928, 83929, 83930, 
    83931, 83932, 83933, 83934, 83935, 83936, 83937, 83938, 83939, 83940, 
    83941, 83942, 83943, 83944, 83945, 83946, 83947, 83948, 83949, 83950, 
    83951, 83952, 83953, 83954, 83955, 83956, 83957, 83958, 83959, 83960, 
    83961, 83962, 83963, 83964, 83965, 83966, 83967, 83968, 83969, 83970, 
    83971, 83972, 83973, 83974, 83975, 83976, 83977, 83978, 83979, 83980, 
    83981, 83982, 83983, 83984, 83985, 83986, 83987, 83988, 83989, 83990, 
    83991, 83992, 83993, 83994, 83995, 83996, 83997, 83998, 83999, 84000, 
    84001, 84002, 84003, 84004, 84005, 84006, 84007, 84008, 84009, 84010, 
    84011, 84012, 84013, 84014, 84015, 84016, 84017, 84018, 84019, 84020, 
    84021, 84022, 84023, 84024, 84025, 84026, 84027, 84028, 84029, 84030, 
    84031, 84032, 84033, 84034, 84035, 84036, 84037, 84038, 84039, 84040, 
    84041, 84042, 84043, 84044, 84045, 84046, 84047, 84048, 84049, 84050, 
    84051, 84052, 84053, 84054, 84055, 84056, 84057, 84058, 84059, 84060, 
    84061, 84062, 84063, 84064, 84065, 84066, 84067, 84068, 84069, 84070, 
    84071, 84072, 84073, 84074, 84075, 84076, 84077, 84078, 84079, 84080, 
    84081, 84082, 84083, 84084, 84085, 84086, 84087, 84088, 84089, 84090, 
    84091, 84092, 84093, 84094, 84095, 84096, 84097, 84098, 84099, 84100, 
    84101, 84102, 84103, 84104, 84105, 84106, 84107, 84108, 84109, 84110, 
    84111, 84112, 84113, 84114, 84115, 84116, 84117, 84118, 84119, 84120, 
    84121, 84122, 84123, 84124, 84125, 84126, 84127, 84128, 84129, 84130, 
    84131, 84132, 84133, 84134, 84135, 84136, 84137, 84138, 84139, 84140, 
    84141, 84142, 84143, 84144, 84145, 84146, 84147, 84148, 84149, 84150, 
    84151, 84152, 84153, 84154, 84155, 84156, 84157, 84158, 84159, 84160, 
    84161, 84162, 84163, 84164, 84165, 84166, 84167, 84168, 84169, 84170, 
    84171, 84172, 84173, 84174, 84175, 84176, 84177, 84178, 84179, 84180, 
    84181, 84182, 84183, 84184, 84185, 84186, 84187, 84188, 84189, 84190, 
    84191, 84192, 84193, 84194, 84195, 84196, 84197, 84198, 84199, 84200, 
    84201, 84202, 84203, 84204, 84205, 84206, 84207, 84208, 84209, 84210, 
    84211, 84212, 84213, 84214, 84215, 84216, 84217, 84218, 84219, 84220, 
    84221, 84222, 84223, 84224, 84225, 84226, 84227, 84228, 84229, 84230, 
    84231, 84232, 84233, 84234, 84235, 84236, 84237, 84238, 84239, 84240, 
    84241, 84242, 84243, 84244, 84245, 84246, 84247, 84248, 84249, 84250, 
    84251, 84252, 84253, 84254, 84255, 84256, 84257, 84258, 84259, 84260, 
    84261, 84262, 84263, 84264, 84265, 84266, 84267, 84268, 84269, 84270, 
    84271, 84272, 84273, 84274, 84275, 84276, 84277, 84278, 84279, 84280, 
    84281, 84282, 84283, 84284, 84285, 84286, 84287, 84288, 84289, 84290, 
    84291, 84292, 84293, 84294, 84295, 84296, 84297, 84298, 84299, 84300, 
    84301, 84302, 84303, 84304, 84305, 84306, 84307, 84308, 84309, 84310, 
    84311, 84312, 84313, 84314, 84315, 84316, 84317, 84318, 84319, 84320, 
    84321, 84322, 84323, 84324, 84325, 84326, 84327, 84328, 84329, 84330, 
    84331, 84332, 84333, 84334, 84335, 84336, 84337, 84338, 84339, 84340, 
    84341, 84342, 84343, 84344, 84345, 84346, 84347, 84348, 84349, 84350, 
    84351, 84352, 84353, 84354, 84355, 84356, 84357, 84358, 84359, 84360, 
    84361, 84362, 84363, 84364, 84365, 84366, 84367, 84368, 84369, 84370, 
    84371, 84372, 84373, 84374, 84375, 84376, 84377, 84378, 84379, 84380, 
    84381, 84382, 84383, 84384, 84385, 84386, 84387, 84388, 84389, 84390, 
    84391, 84392, 84393, 84394, 84395, 84396, 84397, 84398, 84399, 84400, 
    84401, 84402, 84403, 84404, 84405, 84406, 84407, 84408, 84409, 84410, 
    84411, 84412, 84413, 84414, 84415, 84416, 84417, 84418, 84419, 84420, 
    84421, 84422, 84423, 84424, 84425, 84426, 84427, 84428, 84429, 84430, 
    84431, 84432, 84433, 84434, 84435, 84436, 84437, 84438, 84439, 84440, 
    84441, 84442, 84443, 84444, 84445, 84446, 84447, 84448, 84449, 84450, 
    84451, 84452, 84453, 84454, 84455, 84456, 84457, 84458, 84459, 84460, 
    84461, 84462, 84463, 84464, 84465, 84466, 84467, 84468, 84469, 84470, 
    84471, 84472, 84473, 84474, 84475, 84476, 84477, 84478, 84479, 84480, 
    84481, 84482, 84483, 84484, 84485, 84486, 84487, 84488, 84489, 84490, 
    84491, 84492, 84493, 84494, 84495, 84496, 84497, 84498, 84499, 84500, 
    84501, 84502, 84503, 84504, 84505, 84506, 84507, 84508, 84509, 84510, 
    84511, 84512, 84513, 84514, 84515, 84516, 84517, 84518, 84519, 84520, 
    84521, 84522, 84523, 84524, 84525, 84526, 84527, 84528, 84529, 84530, 
    84531, 84532, 84533, 84534, 84535, 84536, 84537, 84538, 84539, 84540, 
    84541, 84542, 84543, 84544, 84545, 84546, 84547, 84548, 84549, 84550, 
    84551, 84552, 84553, 84554, 84555, 84556, 84557, 84558, 84559, 84560, 
    84561, 84562, 84563, 84564, 84565, 84566, 84567, 84568, 84569, 84570, 
    84571, 84572, 84573, 84574, 84575, 84576, 84577, 84578, 84579, 84580, 
    84581, 84582, 84583, 84584, 84585, 84586, 84587, 84588, 84589, 84590, 
    84591, 84592, 84593, 84594, 84595, 84596, 84597, 84598, 84599, 84600, 
    84601, 84602, 84603, 84604, 84605, 84606, 84607, 84608, 84609, 84610, 
    84611, 84612, 84613, 84614, 84615, 84616, 84617, 84618, 84619, 84620, 
    84621, 84622, 84623, 84624, 84625, 84626, 84627, 84628, 84629, 84630, 
    84631, 84632, 84633, 84634, 84635, 84636, 84637, 84638, 84639, 84640, 
    84641, 84642, 84643, 84644, 84645, 84646, 84647, 84648, 84649, 84650, 
    84651, 84652, 84653, 84654, 84655, 84656, 84657, 84658, 84659, 84660, 
    84661, 84662, 84663, 84664, 84665, 84666, 84667, 84668, 84669, 84670, 
    84671, 84672, 84673, 84674, 84675, 84676, 84677, 84678, 84679, 84680, 
    84681, 84682, 84683, 84684, 84685, 84686, 84687, 84688, 84689, 84690, 
    84691, 84692, 84693, 84694, 84695, 84696, 84697, 84698, 84699, 84700, 
    84701, 84702, 84703, 84704, 84705, 84706, 84707, 84708, 84709, 84710, 
    84711, 84712, 84713, 84714, 84715, 84716, 84717, 84718, 84719, 84720, 
    84721, 84722, 84723, 84724, 84725, 84726, 84727, 84728, 84729, 84730, 
    84731, 84732, 84733, 84734, 84735, 84736, 84737, 84738, 84739, 84740, 
    84741, 84742, 84743, 84744, 84745, 84746, 84747, 84748, 84749, 84750, 
    84751, 84752, 84753, 84754, 84755, 84756, 84757, 84758, 84759, 84760, 
    84761, 84762, 84763, 84764, 84765, 84766, 84767, 84768, 84769, 84770, 
    84771, 84772, 84773, 84774, 84775, 84776, 84777, 84778, 84779, 84780, 
    84781, 84782, 84783, 84784, 84785, 84786, 84787, 84788, 84789, 84790, 
    84791, 84792, 84793, 84794, 84795, 84796, 84797, 84798, 84799, 84800, 
    84801, 84802, 84803, 84804, 84805, 84806, 84807, 84808, 84809, 84810, 
    84811, 84812, 84813, 84814, 84815, 84816, 84817, 84818, 84819, 84820, 
    84821, 84822, 84823, 84824, 84825, 84826, 84827, 84828, 84829, 84830, 
    84831, 84832, 84833, 84834, 84835, 84836, 84837, 84838, 84839, 84840, 
    84841, 84842, 84843, 84844, 84845, 84846, 84847, 84848, 84849, 84850, 
    84851, 84852, 84853, 84854, 84855, 84856, 84857, 84858, 84859, 84860, 
    84861, 84862, 84863, 84864, 84865, 84866, 84867, 84868, 84869, 84870, 
    84871, 84872, 84873, 84874, 84875, 84876, 84877, 84878, 84879, 84880, 
    84881, 84882, 84883, 84884, 84885, 84886, 84887, 84888, 84889, 84890, 
    84891, 84892, 84893, 84894, 84895, 84896, 84897, 84898, 84899, 84900, 
    84901, 84902, 84903, 84904, 84905, 84906, 84907, 84908, 84909, 84910, 
    84911, 84912, 84913, 84914, 84915, 84916, 84917, 84918, 84919, 84920, 
    84921, 84922, 84923, 84924, 84925, 84926, 84927, 84928, 84929, 84930, 
    84931, 84932, 84933, 84934, 84935, 84936, 84937, 84938, 84939, 84940, 
    84941, 84942, 84943, 84944, 84945, 84946, 84947, 84948, 84949, 84950, 
    84951, 84952, 84953, 84954, 84955, 84956, 84957, 84958, 84959, 84960, 
    84961, 84962, 84963, 84964, 84965, 84966, 84967, 84968, 84969, 84970, 
    84971, 84972, 84973, 84974, 84975, 84976, 84977, 84978, 84979, 84980, 
    84981, 84982, 84983, 84984, 84985, 84986, 84987, 84988, 84989, 84990, 
    84991, 84992, 84993, 84994, 84995, 84996, 84997, 84998, 84999, 85000, 
    85001, 85002, 85003, 85004, 85005, 85006, 85007, 85008, 85009, 85010, 
    85011, 85012, 85013, 85014, 85015, 85016, 85017, 85018, 85019, 85020, 
    85021, 85022, 85023, 85024, 85025, 85026, 85027, 85028, 85029, 85030, 
    85031, 85032, 85033, 85034, 85035, 85036, 85037, 85038, 85039, 85040, 
    85041, 85042, 85043, 85044, 85045, 85046, 85047, 85048, 85049, 85050, 
    85051, 85052, 85053, 85054, 85055, 85056, 85057, 85058, 85059, 85060, 
    85061, 85062, 85063, 85064, 85065, 85066, 85067, 85068, 85069, 85070, 
    85071, 85072, 85073, 85074, 85075, 85076, 85077, 85078, 85079, 85080, 
    85081, 85082, 85083, 85084, 85085, 85086, 85087, 85088, 85089, 85090, 
    85091, 85092, 85093, 85094, 85095, 85096, 85097, 85098, 85099, 85100, 
    85101, 85102, 85103, 85104, 85105, 85106, 85107, 85108, 85109, 85110, 
    85111, 85112, 85113, 85114, 85115, 85116, 85117, 85118, 85119, 85120, 
    85121, 85122, 85123, 85124, 85125, 85126, 85127, 85128, 85129, 85130, 
    85131, 85132, 85133, 85134, 85135, 85136, 85137, 85138, 85139, 85140, 
    85141, 85142, 85143, 85144, 85145, 85146, 85147, 85148, 85149, 85150, 
    85151, 85152, 85153, 85154, 85155, 85156, 85157, 85158, 85159, 85160, 
    85161, 85162, 85163, 85164, 85165, 85166, 85167, 85168, 85169, 85170, 
    85171, 85172, 85173, 85174, 85175, 85176, 85177, 85178, 85179, 85180, 
    85181, 85182, 85183, 85184, 85185, 85186, 85187, 85188, 85189, 85190, 
    85191, 85192, 85193, 85194, 85195, 85196, 85197, 85198, 85199, 85200, 
    85201, 85202, 85203, 85204, 85205, 85206, 85207, 85208, 85209, 85210, 
    85211, 85212, 85213, 85214, 85215, 85216, 85217, 85218, 85219, 85220, 
    85221, 85222, 85223, 85224, 85225, 85226, 85227, 85228, 85229, 85230, 
    85231, 85232, 85233, 85234, 85235, 85236, 85237, 85238, 85239, 85240, 
    85241, 85242, 85243, 85244, 85245, 85246, 85247, 85248, 85249, 85250, 
    85251, 85252, 85253, 85254, 85255, 85256, 85257, 85258, 85259, 85260, 
    85261, 85262, 85263, 85264, 85265, 85266, 85267, 85268, 85269, 85270, 
    85271, 85272, 85273, 85274, 85275, 85276, 85277, 85278, 85279, 85280, 
    85281, 85282, 85283, 85284, 85285, 85286, 85287, 85288, 85289, 85290, 
    85291, 85292, 85293, 85294, 85295, 85296, 85297, 85298, 85299, 85300, 
    85301, 85302, 85303, 85304, 85305, 85306, 85307, 85308, 85309, 85310, 
    85311, 85312, 85313, 85314, 85315, 85316, 85317, 85318, 85319, 85320, 
    85321, 85322, 85323, 85324, 85325, 85326, 85327, 85328, 85329, 85330, 
    85331, 85332, 85333, 85334, 85335, 85336, 85337, 85338, 85339, 85340, 
    85341, 85342, 85343, 85344, 85345, 85346, 85347, 85348, 85349, 85350, 
    85351, 85352, 85353, 85354, 85355, 85356, 85357, 85358, 85359, 85360, 
    85361, 85362, 85363, 85364, 85365, 85366, 85367, 85368, 85369, 85370, 
    85371, 85372, 85373, 85374, 85375, 85376, 85377, 85378, 85379, 85380, 
    85381, 85382, 85383, 85384, 85385, 85386, 85387, 85388, 85389, 85390, 
    85391, 85392, 85393, 85394, 85395, 85396, 85397, 85398, 85399, 85400, 
    85401, 85402, 85403, 85404, 85405, 85406, 85407, 85408, 85409, 85410, 
    85411, 85412, 85413, 85414, 85415, 85416, 85417, 85418, 85419, 85420, 
    85421, 85422, 85423, 85424, 85425, 85426, 85427, 85428, 85429, 85430, 
    85431, 85432, 85433, 85434, 85435, 85436, 85437, 85438, 85439, 85440, 
    85441, 85442, 85443, 85444, 85445, 85446, 85447, 85448, 85449, 85450, 
    85451, 85452, 85453, 85454, 85455, 85456, 85457, 85458, 85459, 85460, 
    85461, 85462, 85463, 85464, 85465, 85466, 85467, 85468, 85469, 85470, 
    85471, 85472, 85473, 85474, 85475, 85476, 85477, 85478, 85479, 85480, 
    85481, 85482, 85483, 85484, 85485, 85486, 85487, 85488, 85489, 85490, 
    85491, 85492, 85493, 85494, 85495, 85496, 85497, 85498, 85499, 85500, 
    85501, 85502, 85503, 85504, 85505, 85506, 85507, 85508, 85509, 85510, 
    85511, 85512, 85513, 85514, 85515, 85516, 85517, 85518, 85519, 85520, 
    85521, 85522, 85523, 85524, 85525, 85526, 85527, 85528, 85529, 85530, 
    85531, 85532, 85533, 85534, 85535, 85536, 85537, 85538, 85539, 85540, 
    85541, 85542, 85543, 85544, 85545, 85546, 85547, 85548, 85549, 85550, 
    85551, 85552, 85553, 85554, 85555, 85556, 85557, 85558, 85559, 85560, 
    85561, 85562, 85563, 85564, 85565, 85566, 85567, 85568, 85569, 85570, 
    85571, 85572, 85573, 85574, 85575, 85576, 85577, 85578, 85579, 85580, 
    85581, 85582, 85583, 85584, 85585, 85586, 85587, 85588, 85589, 85590, 
    85591, 85592, 85593, 85594, 85595, 85596, 85597, 85598, 85599, 85600, 
    85601, 85602, 85603, 85604, 85605, 85606, 85607, 85608, 85609, 85610, 
    85611, 85612, 85613, 85614, 85615, 85616, 85617, 85618, 85619, 85620, 
    85621, 85622, 85623, 85624, 85625, 85626, 85627, 85628, 85629, 85630, 
    85631, 85632, 85633, 85634, 85635, 85636, 85637, 85638, 85639, 85640, 
    85641, 85642, 85643, 85644, 85645, 85646, 85647, 85648, 85649, 85650, 
    85651, 85652, 85653, 85654, 85655, 85656, 85657, 85658, 85659, 85660, 
    85661, 85662, 85663, 85664, 85665, 85666, 85667, 85668, 85669, 85670, 
    85671, 85672, 85673, 85674, 85675, 85676, 85677, 85678, 85679, 85680, 
    85681, 85682, 85683, 85684, 85685, 85686, 85687, 85688, 85689, 85690, 
    85691, 85692, 85693, 85694, 85695, 85696, 85697, 85698, 85699, 85700, 
    85701, 85702, 85703, 85704, 85705, 85706, 85707, 85708, 85709, 85710, 
    85711, 85712, 85713, 85714, 85715, 85716, 85717, 85718, 85719, 85720, 
    85721, 85722, 85723, 85724, 85725, 85726, 85727, 85728, 85729, 85730, 
    85731, 85732, 85733, 85734, 85735, 85736, 85737, 85738, 85739, 85740, 
    85741, 85742, 85743, 85744, 85745, 85746, 85747, 85748, 85749, 85750, 
    85751, 85752, 85753, 85754, 85755, 85756, 85757, 85758, 85759, 85760, 
    85761, 85762, 85763, 85764, 85765, 85766, 85767, 85768, 85769, 85770, 
    85771, 85772, 85773, 85774, 85775, 85776, 85777, 85778, 85779, 85780, 
    85781, 85782, 85783, 85784, 85785, 85786, 85787, 85788, 85789, 85790, 
    85791, 85792, 85793, 85794, 85795, 85796, 85797, 85798, 85799, 85800, 
    85801, 85802, 85803, 85804, 85805, 85806, 85807, 85808, 85809, 85810, 
    85811, 85812, 85813, 85814, 85815, 85816, 85817, 85818, 85819, 85820, 
    85821, 85822, 85823, 85824, 85825, 85826, 85827, 85828, 85829, 85830, 
    85831, 85832, 85833, 85834, 85835, 85836, 85837, 85838, 85839, 85840, 
    85841, 85842, 85843, 85844, 85845, 85846, 85847, 85848, 85849, 85850, 
    85851, 85852, 85853, 85854, 85855, 85856, 85857, 85858, 85859, 85860, 
    85861, 85862, 85863, 85864, 85865, 85866, 85867, 85868, 85869, 85870, 
    85871, 85872, 85873, 85874, 85875, 85876, 85877, 85878, 85879, 85880, 
    85881, 85882, 85883, 85884, 85885, 85886, 85887, 85888, 85889, 85890, 
    85891, 85892, 85893, 85894, 85895, 85896, 85897, 85898, 85899, 85900, 
    85901, 85902, 85903, 85904, 85905, 85906, 85907, 85908, 85909, 85910, 
    85911, 85912, 85913, 85914, 85915, 85916, 85917, 85918, 85919, 85920, 
    85921, 85922, 85923, 85924, 85925, 85926, 85927, 85928, 85929, 85930, 
    85931, 85932, 85933, 85934, 85935, 85936, 85937, 85938, 85939, 85940, 
    85941, 85942, 85943, 85944, 85945, 85946, 85947, 85948, 85949, 85950, 
    85951, 85952, 85953, 85954, 85955, 85956, 85957, 85958, 85959, 85960, 
    85961, 85962, 85963, 85964, 85965, 85966, 85967, 85968, 85969, 85970, 
    85971, 85972, 85973, 85974, 85975, 85976, 85977, 85978, 85979, 85980, 
    85981, 85982, 85983, 85984, 85985, 85986, 85987, 85988, 85989, 85990, 
    85991, 85992, 85993, 85994, 85995, 85996, 85997, 85998, 85999, 86000, 
    86001, 86002, 86003, 86004, 86005, 86006, 86007, 86008, 86009, 86010, 
    86011, 86012, 86013, 86014, 86015, 86016, 86017, 86018, 86019, 86020, 
    86021, 86022, 86023, 86024, 86025, 86026, 86027, 86028, 86029, 86030, 
    86031, 86032, 86033, 86034, 86035, 86036, 86037, 86038, 86039, 86040, 
    86041, 86042, 86043, 86044, 86045, 86046, 86047, 86048, 86049, 86050, 
    86051, 86052, 86053, 86054, 86055, 86056, 86057, 86058, 86059, 86060, 
    86061, 86062, 86063, 86064, 86065, 86066, 86067, 86068, 86069, 86070, 
    86071, 86072, 86073, 86074, 86075, 86076, 86077, 86078, 86079, 86080, 
    86081, 86082, 86083, 86084, 86085, 86086, 86087, 86088, 86089, 86090, 
    86091, 86092, 86093, 86094, 86095, 86096, 86097, 86098, 86099, 86100, 
    86101, 86102, 86103, 86104, 86105, 86106, 86107, 86108, 86109, 86110, 
    86111, 86112, 86113, 86114, 86115, 86116, 86117, 86118, 86119, 86120, 
    86121, 86122, 86123, 86124, 86125, 86126, 86127, 86128, 86129, 86130, 
    86131, 86132, 86133, 86134, 86135, 86136, 86137, 86138, 86139, 86140, 
    86141, 86142, 86143, 86144, 86145, 86146, 86147, 86148, 86149, 86150, 
    86151, 86152, 86153, 86154, 86155, 86156, 86157, 86158, 86159, 86160, 
    86161, 86162, 86163, 86164, 86165, 86166, 86167, 86168, 86169, 86170, 
    86171, 86172, 86173, 86174, 86175, 86176, 86177, 86178, 86179, 86180, 
    86181, 86182, 86183, 86184, 86185, 86186, 86187, 86188, 86189, 86190, 
    86191, 86192, 86193, 86194, 86195, 86196, 86197, 86198, 86199, 86200, 
    86201, 86202, 86203, 86204, 86205, 86206, 86207, 86208, 86209, 86210, 
    86211, 86212, 86213, 86214, 86215, 86216, 86217, 86218, 86219, 86220, 
    86221, 86222, 86223, 86224, 86225, 86226, 86227, 86228, 86229, 86230, 
    86231, 86232, 86233, 86234, 86235, 86236, 86237, 86238, 86239, 86240, 
    86241, 86242, 86243, 86244, 86245, 86246, 86247, 86248, 86249, 86250, 
    86251, 86252, 86253, 86254, 86255, 86256, 86257, 86258, 86259, 86260, 
    86261, 86262, 86263, 86264, 86265, 86266, 86267, 86268, 86269, 86270, 
    86271, 86272, 86273, 86274, 86275, 86276, 86277, 86278, 86279, 86280, 
    86281, 86282, 86283, 86284, 86285, 86286, 86287, 86288, 86289, 86290, 
    86291, 86292, 86293, 86294, 86295, 86296, 86297, 86298, 86299, 86300, 
    86301, 86302, 86303, 86304, 86305, 86306, 86307, 86308, 86309, 86310, 
    86311, 86312, 86313, 86314, 86315, 86316, 86317, 86318, 86319, 86320, 
    86321, 86322, 86323, 86324, 86325, 86326, 86327, 86328, 86329, 86330, 
    86331, 86332, 86333, 86334, 86335, 86336, 86337, 86338, 86339, 86340, 
    86341, 86342, 86343, 86344, 86345, 86346, 86347, 86348, 86349, 86350, 
    86351, 86352, 86353, 86354, 86355, 86356, 86357, 86358, 86359, 86360, 
    86361, 86362, 86363, 86364, 86365, 86366, 86367, 86368, 86369, 86370, 
    86371, 86372, 86373, 86374, 86375, 86376, 86377, 86378, 86379, 86380, 
    86381, 86382, 86383, 86384, 86385, 86386, 86387, 86388, 86389, 86390, 
    86391, 86392, 86393, 86394, 86395, 86396, 86397, 86398, 86399, 86400, 
    86401, 86402, 86403, 86404, 86405, 86406, 86407, 86408, 86409, 86410, 
    86411, 86412, 86413, 86414, 86415, 86416, 86417, 86418, 86419, 86420, 
    86421, 86422, 86423, 86424, 86425, 86426, 86427, 86428, 86429, 86430, 
    86431, 86432, 86433, 86434, 86435, 86436, 86437, 86438, 86439, 86440, 
    86441, 86442, 86443, 86444, 86445, 86446, 86447, 86448, 86449, 86450, 
    86451, 86452, 86453, 86454, 86455, 86456, 86457, 86458, 86459, 86460, 
    86461, 86462, 86463, 86464, 86465, 86466, 86467, 86468, 86469, 86470, 
    86471, 86472, 86473, 86474, 86475, 86476, 86477, 86478, 86479, 86480, 
    86481, 86482, 86483, 86484, 86485, 86486, 86487, 86488, 86489, 86490, 
    86491, 86492, 86493, 86494, 86495, 86496, 86497, 86498, 86499, 86500, 
    86501, 86502, 86503, 86504, 86505, 86506, 86507, 86508, 86509, 86510, 
    86511, 86512, 86513, 86514, 86515, 86516, 86517, 86518, 86519, 86520, 
    86521, 86522, 86523, 86524, 86525, 86526, 86527, 86528, 86529, 86530, 
    86531, 86532, 86533, 86534, 86535, 86536, 86537, 86538, 86539, 86540, 
    86541, 86542, 86543, 86544, 86545, 86546, 86547, 86548, 86549, 86550, 
    86551, 86552, 86553, 86554, 86555, 86556, 86557, 86558, 86559, 86560, 
    86561, 86562, 86563, 86564, 86565, 86566, 86567, 86568, 86569, 86570, 
    86571, 86572, 86573, 86574, 86575, 86576, 86577, 86578, 86579, 86580, 
    86581, 86582, 86583, 86584, 86585, 86586, 86587, 86588, 86589, 86590, 
    86591, 86592, 86593, 86594, 86595, 86596, 86597, 86598, 86599, 86600, 
    86601, 86602, 86603, 86604, 86605, 86606, 86607, 86608, 86609, 86610, 
    86611, 86612, 86613, 86614, 86615, 86616, 86617, 86618, 86619, 86620, 
    86621, 86622, 86623, 86624, 86625, 86626, 86627, 86628, 86629, 86630, 
    86631, 86632, 86633, 86634, 86635, 86636, 86637, 86638, 86639, 86640, 
    86641, 86642, 86643, 86644, 86645, 86646, 86647, 86648, 86649, 86650, 
    86651, 86652, 86653, 86654, 86655, 86656, 86657, 86658, 86659, 86660, 
    86661, 86662, 86663, 86664, 86665, 86666, 86667, 86668, 86669, 86670, 
    86671, 86672, 86673, 86674, 86675, 86676, 86677, 86678, 86679, 86680, 
    86681, 86682, 86683, 86684, 86685, 86686, 86687, 86688, 86689, 86690, 
    86691, 86692, 86693, 86694, 86695, 86696, 86697, 86698, 86699, 86700, 
    86701, 86702, 86703, 86704, 86705, 86706, 86707, 86708, 86709, 86710, 
    86711, 86712, 86713, 86714, 86715, 86716, 86717, 86718, 86719, 86720, 
    86721, 86722, 86723, 86724, 86725, 86726, 86727, 86728, 86729, 86730, 
    86731, 86732, 86733, 86734, 86735, 86736, 86737, 86738, 86739, 86740, 
    86741, 86742, 86743, 86744, 86745, 86746, 86747, 86748, 86749, 86750, 
    86751, 86752, 86753, 86754, 86755, 86756, 86757, 86758, 86759, 86760, 
    86761, 86762, 86763, 86764, 86765, 86766, 86767, 86768, 86769, 86770, 
    86771, 86772, 86773, 86774, 86775, 86776, 86777, 86778, 86779, 86780, 
    86781, 86782, 86783, 86784, 86785, 86786, 86787, 86788, 86789, 86790, 
    86791, 86792, 86793, 86794, 86795, 86796, 86797, 86798, 86799, 86800, 
    86801, 86802, 86803, 86804, 86805, 86806, 86807, 86808, 86809, 86810, 
    86811, 86812, 86813, 86814, 86815, 86816, 86817, 86818, 86819, 86820, 
    86821, 86822, 86823, 86824, 86825, 86826, 86827, 86828, 86829, 86830, 
    86831, 86832, 86833, 86834, 86835, 86836, 86837, 86838, 86839, 86840, 
    86841, 86842, 86843, 86844, 86845, 86846, 86847, 86848, 86849, 86850, 
    86851, 86852, 86853, 86854, 86855, 86856, 86857, 86858, 86859, 86860, 
    86861, 86862, 86863, 86864, 86865, 86866, 86867, 86868, 86869, 86870, 
    86871, 86872, 86873, 86874, 86875, 86876, 86877, 86878, 86879, 86880, 
    86881, 86882, 86883, 86884, 86885, 86886, 86887, 86888, 86889, 86890, 
    86891, 86892, 86893, 86894, 86895, 86896, 86897, 86898, 86899, 86900, 
    86901, 86902, 86903, 86904, 86905, 86906, 86907, 86908, 86909, 86910, 
    86911, 86912, 86913, 86914, 86915, 86916, 86917, 86918, 86919, 86920, 
    86921, 86922, 86923, 86924, 86925, 86926, 86927, 86928, 86929, 86930, 
    86931, 86932, 86933, 86934, 86935, 86936, 86937, 86938, 86939, 86940, 
    86941, 86942, 86943, 86944, 86945, 86946, 86947, 86948, 86949, 86950, 
    86951, 86952, 86953, 86954, 86955, 86956, 86957, 86958, 86959, 86960, 
    86961, 86962, 86963, 86964, 86965, 86966, 86967, 86968, 86969, 86970, 
    86971, 86972, 86973, 86974, 86975, 86976, 86977, 86978, 86979, 86980, 
    86981, 86982, 86983, 86984, 86985, 86986, 86987, 86988, 86989, 86990, 
    86991, 86992, 86993, 86994, 86995, 86996, 86997, 86998, 86999, 87000, 
    87001, 87002, 87003, 87004, 87005, 87006, 87007, 87008, 87009, 87010, 
    87011, 87012, 87013, 87014, 87015, 87016, 87017, 87018, 87019, 87020, 
    87021, 87022, 87023, 87024, 87025, 87026, 87027, 87028, 87029, 87030, 
    87031, 87032, 87033, 87034, 87035, 87036, 87037, 87038, 87039, 87040, 
    87041, 87042, 87043, 87044, 87045, 87046, 87047, 87048, 87049, 87050, 
    87051, 87052, 87053, 87054, 87055, 87056, 87057, 87058, 87059, 87060, 
    87061, 87062, 87063, 87064, 87065, 87066, 87067, 87068, 87069, 87070, 
    87071, 87072, 87073, 87074, 87075, 87076, 87077, 87078, 87079, 87080, 
    87081, 87082, 87083, 87084, 87085, 87086, 87087, 87088, 87089, 87090, 
    87091, 87092, 87093, 87094, 87095, 87096, 87097, 87098, 87099, 87100, 
    87101, 87102, 87103, 87104, 87105, 87106, 87107, 87108, 87109, 87110, 
    87111, 87112, 87113, 87114, 87115, 87116, 87117, 87118, 87119, 87120, 
    87121, 87122, 87123, 87124, 87125, 87126, 87127, 87128, 87129, 87130, 
    87131, 87132, 87133, 87134, 87135, 87136, 87137, 87138, 87139, 87140, 
    87141, 87142, 87143, 87144, 87145, 87146, 87147, 87148, 87149, 87150, 
    87151, 87152, 87153, 87154, 87155, 87156, 87157, 87158, 87159, 87160, 
    87161, 87162, 87163, 87164, 87165, 87166, 87167, 87168, 87169, 87170, 
    87171, 87172, 87173, 87174, 87175, 87176, 87177, 87178, 87179, 87180, 
    87181, 87182, 87183, 87184, 87185, 87186, 87187, 87188, 87189, 87190, 
    87191, 87192, 87193, 87194, 87195, 87196, 87197, 87198, 87199, 87200, 
    87201, 87202, 87203, 87204, 87205, 87206, 87207, 87208, 87209, 87210, 
    87211, 87212, 87213, 87214, 87215, 87216, 87217, 87218, 87219, 87220, 
    87221, 87222, 87223, 87224, 87225, 87226, 87227, 87228, 87229, 87230, 
    87231, 87232, 87233, 87234, 87235, 87236, 87237, 87238, 87239, 87240, 
    87241, 87242, 87243, 87244, 87245, 87246, 87247, 87248, 87249, 87250, 
    87251, 87252, 87253, 87254, 87255, 87256, 87257, 87258, 87259, 87260, 
    87261, 87262, 87263, 87264, 87265, 87266, 87267, 87268, 87269, 87270, 
    87271, 87272, 87273, 87274, 87275, 87276, 87277, 87278, 87279, 87280, 
    87281, 87282, 87283, 87284, 87285, 87286, 87287, 87288, 87289, 87290, 
    87291, 87292, 87293, 87294, 87295, 87296, 87297, 87298, 87299, 87300, 
    87301, 87302, 87303, 87304, 87305, 87306, 87307, 87308, 87309, 87310, 
    87311, 87312, 87313, 87314, 87315, 87316, 87317, 87318, 87319, 87320, 
    87321, 87322, 87323, 87324, 87325, 87326, 87327, 87328, 87329, 87330, 
    87331, 87332, 87333, 87334, 87335, 87336, 87337, 87338, 87339, 87340, 
    87341, 87342, 87343, 87344, 87345, 87346, 87347, 87348, 87349, 87350, 
    87351, 87352, 87353, 87354, 87355, 87356, 87357, 87358, 87359, 87360, 
    87361, 87362, 87363, 87364, 87365, 87366, 87367, 87368, 87369, 87370, 
    87371, 87372, 87373, 87374, 87375, 87376, 87377, 87378, 87379, 87380, 
    87381, 87382, 87383, 87384, 87385, 87386, 87387, 87388, 87389, 87390, 
    87391, 87392, 87393, 87394, 87395, 87396, 87397, 87398, 87399, 87400, 
    87401, 87402, 87403, 87404, 87405, 87406, 87407, 87408, 87409, 87410, 
    87411, 87412, 87413, 87414, 87415, 87416, 87417, 87418, 87419, 87420, 
    87421, 87422, 87423, 87424, 87425, 87426, 87427, 87428, 87429, 87430, 
    87431, 87432, 87433, 87434, 87435, 87436, 87437, 87438, 87439, 87440, 
    87441, 87442, 87443, 87444, 87445, 87446, 87447, 87448, 87449, 87450, 
    87451, 87452, 87453, 87454, 87455, 87456, 87457, 87458, 87459, 87460, 
    87461, 87462, 87463, 87464, 87465, 87466, 87467, 87468, 87469, 87470, 
    87471, 87472, 87473, 87474, 87475, 87476, 87477, 87478, 87479, 87480, 
    87481, 87482, 87483, 87484, 87485, 87486, 87487, 87488, 87489, 87490, 
    87491, 87492, 87493, 87494, 87495, 87496, 87497, 87498, 87499, 87500, 
    87501, 87502, 87503, 87504, 87505, 87506, 87507, 87508, 87509, 87510, 
    87511, 87512, 87513, 87514, 87515, 87516, 87517, 87518, 87519, 87520, 
    87521, 87522, 87523, 87524, 87525, 87526, 87527, 87528, 87529, 87530, 
    87531, 87532, 87533, 87534, 87535, 87536, 87537, 87538, 87539, 87540, 
    87541, 87542, 87543, 87544, 87545, 87546, 87547, 87548, 87549, 87550, 
    87551, 87552, 87553, 87554, 87555, 87556, 87557, 87558, 87559, 87560, 
    87561, 87562, 87563, 87564, 87565, 87566, 87567, 87568, 87569, 87570, 
    87571, 87572, 87573, 87574, 87575, 87576, 87577, 87578, 87579, 87580, 
    87581, 87582, 87583, 87584, 87585, 87586, 87587, 87588, 87589, 87590, 
    87591, 87592, 87593, 87594, 87595, 87596, 87597, 87598, 87599, 87600, 
    87601, 87602, 87603, 87604, 87605, 87606, 87607, 87608, 87609, 87610, 
    87611, 87612, 87613, 87614, 87615, 87616, 87617, 87618, 87619, 87620, 
    87621, 87622, 87623, 87624, 87625, 87626, 87627, 87628, 87629, 87630, 
    87631, 87632, 87633, 87634, 87635, 87636, 87637, 87638, 87639, 87640, 
    87641, 87642, 87643, 87644, 87645, 87646, 87647, 87648, 87649, 87650, 
    87651, 87652, 87653, 87654, 87655, 87656, 87657, 87658 ;
}
